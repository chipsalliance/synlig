module top(output longint o);
   assign o = 1;
endmodule
