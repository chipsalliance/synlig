module top(output int o);
   import my_pkg::*;
   assign o = A__B;
endmodule
