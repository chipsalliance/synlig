module top(output logic[7:0] o);
   assign o = '{8{1}};
endmodule
