module top(input a, output b);
assign b = a;
endmodule
