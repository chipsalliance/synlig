module top(output int o);
   assign o = 1 + 2;
endmodule
