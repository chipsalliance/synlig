module dut (output logic[63:0] a, output logic[63:0] b, output logic[63:0] c, output logic[63:0] d);
   assign a = 64'd7698294523898761276;
   assign b = 7698294523898761276;
   assign c = 64'b1010110110110101001010101100101010101010101010101010101010101110;
   assign d = 64'hACBF74CFA4B5A09B;
endmodule
