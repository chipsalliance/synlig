module top(input clk, output logic o);
   assign o = logic'(1);
endmodule
