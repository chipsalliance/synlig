module top(output int o);
   always begin
      o = 1;
   end
endmodule // top
