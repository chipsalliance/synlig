

module top
(
  i,
  o
);

  input [15:0] i;
  output [511:0] o;

  bsg_expand_bitmask
  wrapper
  (
    .i(i),
    .o(o)
  );


endmodule



module bsg_expand_bitmask
(
  i,
  o
);

  input [15:0] i;
  output [511:0] o;
  wire [511:0] o;
  wire o_511_,o_479_,o_447_,o_415_,o_383_,o_351_,o_319_,o_287_,o_255_,o_223_,o_191_,
  o_159_,o_127_,o_95_,o_63_,o_31_;
  assign o_511_ = i[15];
  assign o[480] = o_511_;
  assign o[481] = o_511_;
  assign o[482] = o_511_;
  assign o[483] = o_511_;
  assign o[484] = o_511_;
  assign o[485] = o_511_;
  assign o[486] = o_511_;
  assign o[487] = o_511_;
  assign o[488] = o_511_;
  assign o[489] = o_511_;
  assign o[490] = o_511_;
  assign o[491] = o_511_;
  assign o[492] = o_511_;
  assign o[493] = o_511_;
  assign o[494] = o_511_;
  assign o[495] = o_511_;
  assign o[496] = o_511_;
  assign o[497] = o_511_;
  assign o[498] = o_511_;
  assign o[499] = o_511_;
  assign o[500] = o_511_;
  assign o[501] = o_511_;
  assign o[502] = o_511_;
  assign o[503] = o_511_;
  assign o[504] = o_511_;
  assign o[505] = o_511_;
  assign o[506] = o_511_;
  assign o[507] = o_511_;
  assign o[508] = o_511_;
  assign o[509] = o_511_;
  assign o[510] = o_511_;
  assign o[511] = o_511_;
  assign o_479_ = i[14];
  assign o[448] = o_479_;
  assign o[449] = o_479_;
  assign o[450] = o_479_;
  assign o[451] = o_479_;
  assign o[452] = o_479_;
  assign o[453] = o_479_;
  assign o[454] = o_479_;
  assign o[455] = o_479_;
  assign o[456] = o_479_;
  assign o[457] = o_479_;
  assign o[458] = o_479_;
  assign o[459] = o_479_;
  assign o[460] = o_479_;
  assign o[461] = o_479_;
  assign o[462] = o_479_;
  assign o[463] = o_479_;
  assign o[464] = o_479_;
  assign o[465] = o_479_;
  assign o[466] = o_479_;
  assign o[467] = o_479_;
  assign o[468] = o_479_;
  assign o[469] = o_479_;
  assign o[470] = o_479_;
  assign o[471] = o_479_;
  assign o[472] = o_479_;
  assign o[473] = o_479_;
  assign o[474] = o_479_;
  assign o[475] = o_479_;
  assign o[476] = o_479_;
  assign o[477] = o_479_;
  assign o[478] = o_479_;
  assign o[479] = o_479_;
  assign o_447_ = i[13];
  assign o[416] = o_447_;
  assign o[417] = o_447_;
  assign o[418] = o_447_;
  assign o[419] = o_447_;
  assign o[420] = o_447_;
  assign o[421] = o_447_;
  assign o[422] = o_447_;
  assign o[423] = o_447_;
  assign o[424] = o_447_;
  assign o[425] = o_447_;
  assign o[426] = o_447_;
  assign o[427] = o_447_;
  assign o[428] = o_447_;
  assign o[429] = o_447_;
  assign o[430] = o_447_;
  assign o[431] = o_447_;
  assign o[432] = o_447_;
  assign o[433] = o_447_;
  assign o[434] = o_447_;
  assign o[435] = o_447_;
  assign o[436] = o_447_;
  assign o[437] = o_447_;
  assign o[438] = o_447_;
  assign o[439] = o_447_;
  assign o[440] = o_447_;
  assign o[441] = o_447_;
  assign o[442] = o_447_;
  assign o[443] = o_447_;
  assign o[444] = o_447_;
  assign o[445] = o_447_;
  assign o[446] = o_447_;
  assign o[447] = o_447_;
  assign o_415_ = i[12];
  assign o[384] = o_415_;
  assign o[385] = o_415_;
  assign o[386] = o_415_;
  assign o[387] = o_415_;
  assign o[388] = o_415_;
  assign o[389] = o_415_;
  assign o[390] = o_415_;
  assign o[391] = o_415_;
  assign o[392] = o_415_;
  assign o[393] = o_415_;
  assign o[394] = o_415_;
  assign o[395] = o_415_;
  assign o[396] = o_415_;
  assign o[397] = o_415_;
  assign o[398] = o_415_;
  assign o[399] = o_415_;
  assign o[400] = o_415_;
  assign o[401] = o_415_;
  assign o[402] = o_415_;
  assign o[403] = o_415_;
  assign o[404] = o_415_;
  assign o[405] = o_415_;
  assign o[406] = o_415_;
  assign o[407] = o_415_;
  assign o[408] = o_415_;
  assign o[409] = o_415_;
  assign o[410] = o_415_;
  assign o[411] = o_415_;
  assign o[412] = o_415_;
  assign o[413] = o_415_;
  assign o[414] = o_415_;
  assign o[415] = o_415_;
  assign o_383_ = i[11];
  assign o[352] = o_383_;
  assign o[353] = o_383_;
  assign o[354] = o_383_;
  assign o[355] = o_383_;
  assign o[356] = o_383_;
  assign o[357] = o_383_;
  assign o[358] = o_383_;
  assign o[359] = o_383_;
  assign o[360] = o_383_;
  assign o[361] = o_383_;
  assign o[362] = o_383_;
  assign o[363] = o_383_;
  assign o[364] = o_383_;
  assign o[365] = o_383_;
  assign o[366] = o_383_;
  assign o[367] = o_383_;
  assign o[368] = o_383_;
  assign o[369] = o_383_;
  assign o[370] = o_383_;
  assign o[371] = o_383_;
  assign o[372] = o_383_;
  assign o[373] = o_383_;
  assign o[374] = o_383_;
  assign o[375] = o_383_;
  assign o[376] = o_383_;
  assign o[377] = o_383_;
  assign o[378] = o_383_;
  assign o[379] = o_383_;
  assign o[380] = o_383_;
  assign o[381] = o_383_;
  assign o[382] = o_383_;
  assign o[383] = o_383_;
  assign o_351_ = i[10];
  assign o[320] = o_351_;
  assign o[321] = o_351_;
  assign o[322] = o_351_;
  assign o[323] = o_351_;
  assign o[324] = o_351_;
  assign o[325] = o_351_;
  assign o[326] = o_351_;
  assign o[327] = o_351_;
  assign o[328] = o_351_;
  assign o[329] = o_351_;
  assign o[330] = o_351_;
  assign o[331] = o_351_;
  assign o[332] = o_351_;
  assign o[333] = o_351_;
  assign o[334] = o_351_;
  assign o[335] = o_351_;
  assign o[336] = o_351_;
  assign o[337] = o_351_;
  assign o[338] = o_351_;
  assign o[339] = o_351_;
  assign o[340] = o_351_;
  assign o[341] = o_351_;
  assign o[342] = o_351_;
  assign o[343] = o_351_;
  assign o[344] = o_351_;
  assign o[345] = o_351_;
  assign o[346] = o_351_;
  assign o[347] = o_351_;
  assign o[348] = o_351_;
  assign o[349] = o_351_;
  assign o[350] = o_351_;
  assign o[351] = o_351_;
  assign o_319_ = i[9];
  assign o[288] = o_319_;
  assign o[289] = o_319_;
  assign o[290] = o_319_;
  assign o[291] = o_319_;
  assign o[292] = o_319_;
  assign o[293] = o_319_;
  assign o[294] = o_319_;
  assign o[295] = o_319_;
  assign o[296] = o_319_;
  assign o[297] = o_319_;
  assign o[298] = o_319_;
  assign o[299] = o_319_;
  assign o[300] = o_319_;
  assign o[301] = o_319_;
  assign o[302] = o_319_;
  assign o[303] = o_319_;
  assign o[304] = o_319_;
  assign o[305] = o_319_;
  assign o[306] = o_319_;
  assign o[307] = o_319_;
  assign o[308] = o_319_;
  assign o[309] = o_319_;
  assign o[310] = o_319_;
  assign o[311] = o_319_;
  assign o[312] = o_319_;
  assign o[313] = o_319_;
  assign o[314] = o_319_;
  assign o[315] = o_319_;
  assign o[316] = o_319_;
  assign o[317] = o_319_;
  assign o[318] = o_319_;
  assign o[319] = o_319_;
  assign o_287_ = i[8];
  assign o[256] = o_287_;
  assign o[257] = o_287_;
  assign o[258] = o_287_;
  assign o[259] = o_287_;
  assign o[260] = o_287_;
  assign o[261] = o_287_;
  assign o[262] = o_287_;
  assign o[263] = o_287_;
  assign o[264] = o_287_;
  assign o[265] = o_287_;
  assign o[266] = o_287_;
  assign o[267] = o_287_;
  assign o[268] = o_287_;
  assign o[269] = o_287_;
  assign o[270] = o_287_;
  assign o[271] = o_287_;
  assign o[272] = o_287_;
  assign o[273] = o_287_;
  assign o[274] = o_287_;
  assign o[275] = o_287_;
  assign o[276] = o_287_;
  assign o[277] = o_287_;
  assign o[278] = o_287_;
  assign o[279] = o_287_;
  assign o[280] = o_287_;
  assign o[281] = o_287_;
  assign o[282] = o_287_;
  assign o[283] = o_287_;
  assign o[284] = o_287_;
  assign o[285] = o_287_;
  assign o[286] = o_287_;
  assign o[287] = o_287_;
  assign o_255_ = i[7];
  assign o[224] = o_255_;
  assign o[225] = o_255_;
  assign o[226] = o_255_;
  assign o[227] = o_255_;
  assign o[228] = o_255_;
  assign o[229] = o_255_;
  assign o[230] = o_255_;
  assign o[231] = o_255_;
  assign o[232] = o_255_;
  assign o[233] = o_255_;
  assign o[234] = o_255_;
  assign o[235] = o_255_;
  assign o[236] = o_255_;
  assign o[237] = o_255_;
  assign o[238] = o_255_;
  assign o[239] = o_255_;
  assign o[240] = o_255_;
  assign o[241] = o_255_;
  assign o[242] = o_255_;
  assign o[243] = o_255_;
  assign o[244] = o_255_;
  assign o[245] = o_255_;
  assign o[246] = o_255_;
  assign o[247] = o_255_;
  assign o[248] = o_255_;
  assign o[249] = o_255_;
  assign o[250] = o_255_;
  assign o[251] = o_255_;
  assign o[252] = o_255_;
  assign o[253] = o_255_;
  assign o[254] = o_255_;
  assign o[255] = o_255_;
  assign o_223_ = i[6];
  assign o[192] = o_223_;
  assign o[193] = o_223_;
  assign o[194] = o_223_;
  assign o[195] = o_223_;
  assign o[196] = o_223_;
  assign o[197] = o_223_;
  assign o[198] = o_223_;
  assign o[199] = o_223_;
  assign o[200] = o_223_;
  assign o[201] = o_223_;
  assign o[202] = o_223_;
  assign o[203] = o_223_;
  assign o[204] = o_223_;
  assign o[205] = o_223_;
  assign o[206] = o_223_;
  assign o[207] = o_223_;
  assign o[208] = o_223_;
  assign o[209] = o_223_;
  assign o[210] = o_223_;
  assign o[211] = o_223_;
  assign o[212] = o_223_;
  assign o[213] = o_223_;
  assign o[214] = o_223_;
  assign o[215] = o_223_;
  assign o[216] = o_223_;
  assign o[217] = o_223_;
  assign o[218] = o_223_;
  assign o[219] = o_223_;
  assign o[220] = o_223_;
  assign o[221] = o_223_;
  assign o[222] = o_223_;
  assign o[223] = o_223_;
  assign o_191_ = i[5];
  assign o[160] = o_191_;
  assign o[161] = o_191_;
  assign o[162] = o_191_;
  assign o[163] = o_191_;
  assign o[164] = o_191_;
  assign o[165] = o_191_;
  assign o[166] = o_191_;
  assign o[167] = o_191_;
  assign o[168] = o_191_;
  assign o[169] = o_191_;
  assign o[170] = o_191_;
  assign o[171] = o_191_;
  assign o[172] = o_191_;
  assign o[173] = o_191_;
  assign o[174] = o_191_;
  assign o[175] = o_191_;
  assign o[176] = o_191_;
  assign o[177] = o_191_;
  assign o[178] = o_191_;
  assign o[179] = o_191_;
  assign o[180] = o_191_;
  assign o[181] = o_191_;
  assign o[182] = o_191_;
  assign o[183] = o_191_;
  assign o[184] = o_191_;
  assign o[185] = o_191_;
  assign o[186] = o_191_;
  assign o[187] = o_191_;
  assign o[188] = o_191_;
  assign o[189] = o_191_;
  assign o[190] = o_191_;
  assign o[191] = o_191_;
  assign o_159_ = i[4];
  assign o[128] = o_159_;
  assign o[129] = o_159_;
  assign o[130] = o_159_;
  assign o[131] = o_159_;
  assign o[132] = o_159_;
  assign o[133] = o_159_;
  assign o[134] = o_159_;
  assign o[135] = o_159_;
  assign o[136] = o_159_;
  assign o[137] = o_159_;
  assign o[138] = o_159_;
  assign o[139] = o_159_;
  assign o[140] = o_159_;
  assign o[141] = o_159_;
  assign o[142] = o_159_;
  assign o[143] = o_159_;
  assign o[144] = o_159_;
  assign o[145] = o_159_;
  assign o[146] = o_159_;
  assign o[147] = o_159_;
  assign o[148] = o_159_;
  assign o[149] = o_159_;
  assign o[150] = o_159_;
  assign o[151] = o_159_;
  assign o[152] = o_159_;
  assign o[153] = o_159_;
  assign o[154] = o_159_;
  assign o[155] = o_159_;
  assign o[156] = o_159_;
  assign o[157] = o_159_;
  assign o[158] = o_159_;
  assign o[159] = o_159_;
  assign o_127_ = i[3];
  assign o[96] = o_127_;
  assign o[97] = o_127_;
  assign o[98] = o_127_;
  assign o[99] = o_127_;
  assign o[100] = o_127_;
  assign o[101] = o_127_;
  assign o[102] = o_127_;
  assign o[103] = o_127_;
  assign o[104] = o_127_;
  assign o[105] = o_127_;
  assign o[106] = o_127_;
  assign o[107] = o_127_;
  assign o[108] = o_127_;
  assign o[109] = o_127_;
  assign o[110] = o_127_;
  assign o[111] = o_127_;
  assign o[112] = o_127_;
  assign o[113] = o_127_;
  assign o[114] = o_127_;
  assign o[115] = o_127_;
  assign o[116] = o_127_;
  assign o[117] = o_127_;
  assign o[118] = o_127_;
  assign o[119] = o_127_;
  assign o[120] = o_127_;
  assign o[121] = o_127_;
  assign o[122] = o_127_;
  assign o[123] = o_127_;
  assign o[124] = o_127_;
  assign o[125] = o_127_;
  assign o[126] = o_127_;
  assign o[127] = o_127_;
  assign o_95_ = i[2];
  assign o[64] = o_95_;
  assign o[65] = o_95_;
  assign o[66] = o_95_;
  assign o[67] = o_95_;
  assign o[68] = o_95_;
  assign o[69] = o_95_;
  assign o[70] = o_95_;
  assign o[71] = o_95_;
  assign o[72] = o_95_;
  assign o[73] = o_95_;
  assign o[74] = o_95_;
  assign o[75] = o_95_;
  assign o[76] = o_95_;
  assign o[77] = o_95_;
  assign o[78] = o_95_;
  assign o[79] = o_95_;
  assign o[80] = o_95_;
  assign o[81] = o_95_;
  assign o[82] = o_95_;
  assign o[83] = o_95_;
  assign o[84] = o_95_;
  assign o[85] = o_95_;
  assign o[86] = o_95_;
  assign o[87] = o_95_;
  assign o[88] = o_95_;
  assign o[89] = o_95_;
  assign o[90] = o_95_;
  assign o[91] = o_95_;
  assign o[92] = o_95_;
  assign o[93] = o_95_;
  assign o[94] = o_95_;
  assign o[95] = o_95_;
  assign o_63_ = i[1];
  assign o[32] = o_63_;
  assign o[33] = o_63_;
  assign o[34] = o_63_;
  assign o[35] = o_63_;
  assign o[36] = o_63_;
  assign o[37] = o_63_;
  assign o[38] = o_63_;
  assign o[39] = o_63_;
  assign o[40] = o_63_;
  assign o[41] = o_63_;
  assign o[42] = o_63_;
  assign o[43] = o_63_;
  assign o[44] = o_63_;
  assign o[45] = o_63_;
  assign o[46] = o_63_;
  assign o[47] = o_63_;
  assign o[48] = o_63_;
  assign o[49] = o_63_;
  assign o[50] = o_63_;
  assign o[51] = o_63_;
  assign o[52] = o_63_;
  assign o[53] = o_63_;
  assign o[54] = o_63_;
  assign o[55] = o_63_;
  assign o[56] = o_63_;
  assign o[57] = o_63_;
  assign o[58] = o_63_;
  assign o[59] = o_63_;
  assign o[60] = o_63_;
  assign o[61] = o_63_;
  assign o[62] = o_63_;
  assign o[63] = o_63_;
  assign o_31_ = i[0];
  assign o[0] = o_31_;
  assign o[1] = o_31_;
  assign o[2] = o_31_;
  assign o[3] = o_31_;
  assign o[4] = o_31_;
  assign o[5] = o_31_;
  assign o[6] = o_31_;
  assign o[7] = o_31_;
  assign o[8] = o_31_;
  assign o[9] = o_31_;
  assign o[10] = o_31_;
  assign o[11] = o_31_;
  assign o[12] = o_31_;
  assign o[13] = o_31_;
  assign o[14] = o_31_;
  assign o[15] = o_31_;
  assign o[16] = o_31_;
  assign o[17] = o_31_;
  assign o[18] = o_31_;
  assign o[19] = o_31_;
  assign o[20] = o_31_;
  assign o[21] = o_31_;
  assign o[22] = o_31_;
  assign o[23] = o_31_;
  assign o[24] = o_31_;
  assign o[25] = o_31_;
  assign o[26] = o_31_;
  assign o[27] = o_31_;
  assign o[28] = o_31_;
  assign o[29] = o_31_;
  assign o[30] = o_31_;
  assign o[31] = o_31_;

endmodule

