module top;
   initial begin
      $display("Bin number 10 should be printed: %b", 2'd2);
   end
endmodule
