

module top
(
  clk_i,
  reset_i,
  grants_en_i,
  reqs_i,
  grants_o,
  sel_one_hot_o,
  v_o,
  tag_o,
  yumi_i
);

  input [15:0] reqs_i;
  output [15:0] grants_o;
  output [15:0] sel_one_hot_o;
  output [3:0] tag_o;
  input clk_i;
  input reset_i;
  input grants_en_i;
  input yumi_i;
  output v_o;

  bsg_round_robin_arb
  wrapper
  (
    .reqs_i(reqs_i),
    .grants_o(grants_o),
    .sel_one_hot_o(sel_one_hot_o),
    .tag_o(tag_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .grants_en_i(grants_en_i),
    .yumi_i(yumi_i),
    .v_o(v_o)
  );


endmodule



module bsg_round_robin_arb
(
  clk_i,
  reset_i,
  grants_en_i,
  reqs_i,
  grants_o,
  sel_one_hot_o,
  v_o,
  tag_o,
  yumi_i
);

  input [15:0] reqs_i;
  output [15:0] grants_o;
  output [15:0] sel_one_hot_o;
  output [3:0] tag_o;
  input clk_i;
  input reset_i;
  input grants_en_i;
  input yumi_i;
  output v_o;
  wire [15:0] grants_o,sel_one_hot_o;
  wire [3:0] tag_o,last_r;
  wire v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,
  N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,
  N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,
  N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,
  N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,
  N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,
  N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
  N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,
  N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,
  N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,
  N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,
  N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,
  N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,
  N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,
  N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,
  N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,
  N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,
  N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,
  N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,
  N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,
  N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,
  N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,
  N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,
  N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,
  N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,
  N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,
  N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,
  N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,
  N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,
  N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,
  N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,
  N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,
  N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,
  N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,
  N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,
  N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,
  N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,
  N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,
  N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,
  N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,
  N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,
  N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,
  N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,
  N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,
  N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,
  N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,
  N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,
  N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,
  N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,
  N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,
  N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,
  N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,
  N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,
  N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,
  N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,
  N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,
  N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,
  N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,
  N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,
  N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,
  N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,
  N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,
  N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,
  N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,
  N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,
  N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,
  N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,
  N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,
  N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,
  N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,
  N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,
  N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,
  N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
  N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,
  N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,
  N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,
  N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,
  N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,
  N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,
  N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,
  N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,
  N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,
  N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,
  N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,
  N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,
  N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,
  N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,
  N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,
  N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,
  N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,
  N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,
  N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,
  N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,
  N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,
  N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,
  N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,
  N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,
  N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,
  N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,
  N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,
  N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,
  N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,
  N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,
  N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,
  N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,
  N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,
  N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,
  N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,
  N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,
  N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,
  N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,
  N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,
  N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,
  N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,
  N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,
  N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,
  N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,
  N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,
  N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,
  N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
  N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,
  N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,
  N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,
  N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,
  N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,
  N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,
  N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,
  N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,
  N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,
  N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,
  N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,
  N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,
  N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,
  N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,
  N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,
  N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,
  N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,
  N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,
  N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,
  N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,
  N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,
  N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,
  N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,
  N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,
  N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,
  N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,
  N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,
  N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,
  N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,
  N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,N2409,N2410,
  N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422,N2423,
  N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,
  N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,N2449,N2450,
  N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462,N2463,
  N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476,
  N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,N2489,N2490,
  N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502,N2503,
  N2504,N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,
  N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,N2530;
  reg last_r_3_sv2v_reg,last_r_2_sv2v_reg,last_r_1_sv2v_reg,last_r_0_sv2v_reg;
  assign last_r[3] = last_r_3_sv2v_reg;
  assign last_r[2] = last_r_2_sv2v_reg;
  assign last_r[1] = last_r_1_sv2v_reg;
  assign last_r[0] = last_r_0_sv2v_reg;
  assign N261 = N918 & N258;
  assign N262 = N259 & N260;
  assign N263 = N290 & N304;
  assign N264 = N278 & N560;
  assign N265 = N261 & N262;
  assign N266 = N263 & N264;
  assign N267 = N748 & N749;
  assign N268 = N265 & N266;
  assign N269 = N267 & N268;
  assign N274 = N270 & N271;
  assign N275 = N272 & N273;
  assign N276 = N274 & N275;
  assign N277 = N276 & reqs_i[1];
  assign N279 = N270 & N271;
  assign N280 = N272 & N273;
  assign N281 = reqs_i[2] & N278;
  assign N282 = N279 & N280;
  assign N283 = N282 & N281;
  assign N284 = N270 & N271;
  assign N285 = N272 & N273;
  assign N286 = reqs_i[3] & N304;
  assign N287 = N284 & N285;
  assign N288 = N286 & N278;
  assign N289 = N287 & N288;
  assign N291 = N270 & N271;
  assign N292 = N272 & N273;
  assign N293 = reqs_i[4] & N290;
  assign N294 = N291 & N292;
  assign N295 = N293 & N309;
  assign N296 = N294 & N295;
  assign N297 = N270 & N271;
  assign N298 = N272 & N273;
  assign N299 = reqs_i[5] & N260;
  assign N300 = N297 & N298;
  assign N301 = N299 & N263;
  assign N302 = N300 & N301;
  assign N303 = N302 & N278;
  assign N305 = N270 & N271;
  assign N306 = N272 & N273;
  assign N307 = reqs_i[6] & N259;
  assign N308 = N260 & N290;
  assign N309 = N304 & N278;
  assign N310 = N305 & N306;
  assign N311 = N307 & N308;
  assign N312 = N310 & N311;
  assign N313 = N312 & N309;
  assign N314 = N270 & N271;
  assign N315 = N272 & N273;
  assign N316 = N314 & N315;
  assign N317 = N409 & N278;
  assign N318 = N316 & N595;
  assign N319 = N318 & N317;
  assign N320 = N270 & N271;
  assign N321 = N272 & N273;
  assign N322 = N320 & N321;
  assign N323 = N506 & N359;
  assign N324 = N322 & N696;
  assign N325 = N324 & N323;
  assign N326 = N270 & N271;
  assign N327 = N272 & N273;
  assign N328 = N326 & N327;
  assign N329 = N328 & N810;
  assign N330 = N422 & N278;
  assign N331 = N329 & N330;
  assign N332 = N270 & N271;
  assign N333 = N272 & N273;
  assign N334 = N332 & N333;
  assign N335 = N334 & N916;
  assign N336 = N519 & N359;
  assign N337 = N335 & N336;
  assign N338 = N270 & N271;
  assign N339 = N272 & N273;
  assign N340 = N338 & N339;
  assign N341 = N409 & N278;
  assign N342 = N340 & N1027;
  assign N343 = N617 & N341;
  assign N344 = N342 & N343;
  assign N345 = N270 & N271;
  assign N346 = N272 & N273;
  assign N347 = N345 & N346;
  assign N348 = N347 & N1127;
  assign N349 = N718 & N323;
  assign N350 = N348 & N349;
  assign N351 = N270 & N271;
  assign N352 = N272 & N273;
  assign N353 = N351 & N352;
  assign N354 = N353 & N1242;
  assign N355 = N354 & N447;
  assign N356 = N355 & N278;
  assign N357 = N270 & N271;
  assign N358 = N272 & N273;
  assign N359 = N304 & N278;
  assign N360 = N357 & N358;
  assign N361 = N360 & N1349;
  assign N362 = N361 & N544;
  assign N363 = N362 & N359;
  assign N364 = last_r[3] | last_r[2];
  assign N365 = last_r[1] | last_r[0];
  assign N366 = N364 | N365;
  assign N367 = N457 | reqs_i[1];
  assign N368 = N366 | N643;
  assign N369 = N368 | N646;
  assign N370 = N369 | N367;
  assign N372 = last_r[3] | last_r[2];
  assign N373 = last_r[1] | last_r[0];
  assign N374 = reqs_i[15] | reqs_i[14];
  assign N375 = reqs_i[1] | N560;
  assign N376 = N372 | N373;
  assign N377 = N374 | N1464;
  assign N378 = N457 | N375;
  assign N379 = N376 | N377;
  assign N380 = N379 | N646;
  assign N381 = N380 | N378;
  assign N383 = N270 & N271;
  assign N384 = N272 & last_r[0];
  assign N385 = N383 & N384;
  assign N386 = N385 & reqs_i[2];
  assign N387 = N270 & N271;
  assign N388 = N272 & last_r[0];
  assign N389 = reqs_i[3] & N304;
  assign N390 = N387 & N388;
  assign N391 = N390 & N389;
  assign N392 = N270 & N271;
  assign N393 = N272 & last_r[0];
  assign N394 = N392 & N393;
  assign N395 = N486 & N304;
  assign N396 = N394 & N395;
  assign N397 = N270 & N271;
  assign N398 = N272 & last_r[0];
  assign N399 = N397 & N398;
  assign N400 = N584 & N409;
  assign N401 = N399 & N400;
  assign N402 = N270 & N271;
  assign N403 = N272 & last_r[0];
  assign N404 = N402 & N403;
  assign N405 = N404 & N497;
  assign N406 = N405 & N304;
  assign N407 = N270 & N271;
  assign N408 = N272 & last_r[0];
  assign N409 = N290 & N304;
  assign N410 = N407 & N408;
  assign N411 = N410 & N595;
  assign N412 = N411 & N409;
  assign N413 = N270 & N271;
  assign N414 = N272 & last_r[0];
  assign N415 = N413 & N414;
  assign N416 = N506 & N304;
  assign N417 = N415 & N696;
  assign N418 = N417 & N416;
  assign N419 = N270 & N271;
  assign N420 = N272 & last_r[0];
  assign N421 = N419 & N420;
  assign N422 = N604 & N409;
  assign N423 = N421 & N810;
  assign N424 = N423 & N422;
  assign N425 = N270 & N271;
  assign N426 = N272 & last_r[0];
  assign N427 = N425 & N426;
  assign N428 = N427 & N916;
  assign N429 = N519 & N304;
  assign N430 = N428 & N429;
  assign N431 = N270 & N271;
  assign N432 = N272 & last_r[0];
  assign N433 = N431 & N432;
  assign N434 = N433 & N1027;
  assign N435 = N617 & N409;
  assign N436 = N434 & N435;
  assign N437 = N270 & N271;
  assign N438 = N272 & last_r[0];
  assign N439 = N437 & N438;
  assign N440 = N439 & N1127;
  assign N441 = N718 & N416;
  assign N442 = N440 & N441;
  assign N443 = N270 & N271;
  assign N444 = N272 & last_r[0];
  assign N445 = N443 & N444;
  assign N446 = N445 & N1242;
  assign N447 = N832 & N422;
  assign N448 = N446 & N447;
  assign N449 = N270 & N271;
  assign N450 = N272 & last_r[0];
  assign N451 = N449 & N450;
  assign N452 = N451 & N1349;
  assign N453 = N452 & N544;
  assign N454 = N453 & N304;
  assign N455 = last_r[3] | last_r[2];
  assign N456 = last_r[1] | N273;
  assign N457 = reqs_i[3] | reqs_i[2];
  assign N458 = N455 | N456;
  assign N459 = N458 | N643;
  assign N460 = N459 | N646;
  assign N461 = N460 | N457;
  assign N463 = N270 & N271;
  assign N464 = N272 & last_r[0];
  assign N465 = N463 & N464;
  assign N466 = N409 & reqs_i[0];
  assign N467 = N465 & N748;
  assign N468 = N749 & N617;
  assign N469 = N467 & N468;
  assign N470 = N469 & N466;
  assign N471 = last_r[3] | last_r[2];
  assign N472 = last_r[1] | N273;
  assign N473 = N278 | reqs_i[0];
  assign N474 = N471 | N472;
  assign N475 = N457 | N473;
  assign N476 = N474 | N377;
  assign N477 = N476 | N646;
  assign N478 = N477 | N475;
  assign N480 = N270 & N271;
  assign N481 = last_r[1] & N273;
  assign N482 = N480 & N481;
  assign N483 = N482 & reqs_i[3];
  assign N484 = N270 & N271;
  assign N485 = last_r[1] & N273;
  assign N486 = reqs_i[4] & N290;
  assign N487 = N484 & N485;
  assign N488 = N487 & N486;
  assign N489 = N270 & N271;
  assign N490 = last_r[1] & N273;
  assign N491 = N489 & N490;
  assign N492 = N584 & N290;
  assign N493 = N491 & N492;
  assign N494 = N270 & N271;
  assign N495 = last_r[1] & N273;
  assign N496 = N494 & N495;
  assign N497 = N685 & N506;
  assign N498 = N496 & N497;
  assign N499 = N270 & N271;
  assign N500 = last_r[1] & N273;
  assign N501 = N499 & N500;
  assign N502 = N501 & N595;
  assign N503 = N502 & N290;
  assign N504 = N270 & N271;
  assign N505 = last_r[1] & N273;
  assign N506 = N260 & N290;
  assign N507 = N504 & N505;
  assign N508 = N507 & N696;
  assign N509 = N508 & N506;
  assign N510 = N270 & N271;
  assign N511 = last_r[1] & N273;
  assign N512 = N510 & N511;
  assign N513 = N604 & N290;
  assign N514 = N512 & N810;
  assign N515 = N514 & N513;
  assign N516 = N270 & N271;
  assign N517 = last_r[1] & N273;
  assign N518 = N516 & N517;
  assign N519 = N705 & N506;
  assign N520 = N518 & N916;
  assign N521 = N520 & N519;
  assign N522 = N270 & N271;
  assign N523 = last_r[1] & N273;
  assign N524 = N522 & N523;
  assign N525 = N524 & N1027;
  assign N526 = N617 & N290;
  assign N527 = N525 & N526;
  assign N528 = N270 & N271;
  assign N529 = last_r[1] & N273;
  assign N530 = N528 & N529;
  assign N531 = N530 & N1127;
  assign N532 = N718 & N506;
  assign N533 = N531 & N532;
  assign N534 = N270 & N271;
  assign N535 = last_r[1] & N273;
  assign N536 = N534 & N535;
  assign N537 = N536 & N1242;
  assign N538 = N832 & N513;
  assign N539 = N537 & N538;
  assign N540 = N270 & N271;
  assign N541 = last_r[1] & N273;
  assign N542 = N540 & N541;
  assign N543 = N542 & N1349;
  assign N544 = N939 & N519;
  assign N545 = N543 & N544;
  assign N546 = last_r[3] | last_r[2];
  assign N547 = N272 | last_r[0];
  assign N548 = N546 | N547;
  assign N549 = N548 | N643;
  assign N550 = N549 | N646;
  assign N551 = N550 | reqs_i[3];
  assign N553 = N270 & N271;
  assign N554 = last_r[1] & N273;
  assign N555 = N290 & reqs_i[0];
  assign N556 = N553 & N554;
  assign N557 = N556 & N748;
  assign N558 = N557 & N468;
  assign N559 = N558 & N555;
  assign N561 = N270 & N271;
  assign N562 = last_r[1] & N273;
  assign N563 = N290 & reqs_i[1];
  assign N564 = N561 & N562;
  assign N565 = N563 & N560;
  assign N566 = N564 & N748;
  assign N567 = N566 & N468;
  assign N568 = N567 & N565;
  assign N569 = last_r[3] | last_r[2];
  assign N570 = N272 | last_r[0];
  assign N571 = reqs_i[3] | N304;
  assign N572 = N569 | N570;
  assign N573 = N571 | N1951;
  assign N574 = N572 | N377;
  assign N575 = N574 | N646;
  assign N576 = N575 | N573;
  assign N578 = N270 & N271;
  assign N579 = last_r[1] & last_r[0];
  assign N580 = N578 & N579;
  assign N581 = N580 & reqs_i[4];
  assign N582 = N270 & N271;
  assign N583 = last_r[1] & last_r[0];
  assign N584 = reqs_i[5] & N260;
  assign N585 = N582 & N583;
  assign N586 = N585 & N584;
  assign N587 = N270 & N271;
  assign N588 = last_r[1] & last_r[0];
  assign N589 = N587 & N588;
  assign N590 = N685 & N260;
  assign N591 = N589 & N590;
  assign N592 = N270 & N271;
  assign N593 = last_r[1] & last_r[0];
  assign N594 = N592 & N593;
  assign N595 = N799 & N604;
  assign N596 = N594 & N595;
  assign N597 = N270 & N271;
  assign N598 = last_r[1] & last_r[0];
  assign N599 = N597 & N598;
  assign N600 = N599 & N696;
  assign N601 = N600 & N260;
  assign N602 = N270 & N271;
  assign N603 = last_r[1] & last_r[0];
  assign N604 = N259 & N260;
  assign N605 = N602 & N603;
  assign N606 = N605 & N810;
  assign N607 = N606 & N604;
  assign N608 = N270 & N271;
  assign N609 = last_r[1] & last_r[0];
  assign N610 = N608 & N609;
  assign N611 = N705 & N260;
  assign N612 = N610 & N916;
  assign N613 = N612 & N611;
  assign N614 = N270 & N271;
  assign N615 = last_r[1] & last_r[0];
  assign N616 = N614 & N615;
  assign N617 = N819 & N604;
  assign N618 = N616 & N1027;
  assign N619 = N618 & N617;
  assign N620 = N270 & N271;
  assign N621 = last_r[1] & last_r[0];
  assign N622 = N620 & N621;
  assign N623 = N622 & N1127;
  assign N624 = N718 & N260;
  assign N625 = N623 & N624;
  assign N626 = N270 & N271;
  assign N627 = last_r[1] & last_r[0];
  assign N628 = N626 & N627;
  assign N629 = N628 & N1242;
  assign N630 = N832 & N604;
  assign N631 = N629 & N630;
  assign N632 = N270 & N271;
  assign N633 = last_r[1] & last_r[0];
  assign N634 = N632 & N633;
  assign N635 = N634 & N1349;
  assign N636 = N939 & N611;
  assign N637 = N635 & N636;
  assign N638 = last_r[3] | last_r[2];
  assign N639 = N272 | N273;
  assign N640 = N741 | reqs_i[14];
  assign N641 = reqs_i[5] | reqs_i[4];
  assign N642 = N638 | N639;
  assign N643 = N640 | N1464;
  assign N644 = N843 | N641;
  assign N645 = N642 | N643;
  assign N646 = N1051 | N644;
  assign N647 = N645 | N646;
  assign N649 = N270 & N271;
  assign N650 = last_r[1] & last_r[0];
  assign N651 = N649 & N650;
  assign N652 = N651 & N748;
  assign N653 = N652 & N468;
  assign N654 = N653 & reqs_i[0];
  assign N655 = N270 & N271;
  assign N656 = last_r[1] & last_r[0];
  assign N657 = reqs_i[1] & N560;
  assign N658 = N655 & N656;
  assign N659 = N658 & N748;
  assign N660 = N659 & N468;
  assign N661 = N660 & N657;
  assign N662 = N270 & N271;
  assign N663 = last_r[1] & last_r[0];
  assign N664 = reqs_i[2] & N278;
  assign N665 = N662 & N663;
  assign N666 = N664 & N560;
  assign N667 = N665 & N748;
  assign N668 = N667 & N468;
  assign N669 = N668 & N666;
  assign N670 = last_r[3] | last_r[2];
  assign N671 = N272 | N273;
  assign N672 = N290 | reqs_i[2];
  assign N673 = N670 | N671;
  assign N674 = N672 | N1951;
  assign N675 = N673 | N377;
  assign N676 = N675 | N646;
  assign N677 = N676 | N674;
  assign N679 = N270 & last_r[2];
  assign N680 = N272 & N273;
  assign N681 = N679 & N680;
  assign N682 = N681 & reqs_i[5];
  assign N683 = N270 & last_r[2];
  assign N684 = N272 & N273;
  assign N685 = reqs_i[6] & N259;
  assign N686 = N683 & N684;
  assign N687 = N686 & N685;
  assign N688 = N270 & last_r[2];
  assign N689 = N272 & N273;
  assign N690 = N688 & N689;
  assign N691 = N799 & N259;
  assign N692 = N690 & N691;
  assign N693 = N270 & last_r[2];
  assign N694 = N272 & N273;
  assign N695 = N693 & N694;
  assign N696 = N905 & N705;
  assign N697 = N695 & N696;
  assign N698 = N270 & last_r[2];
  assign N699 = N272 & N273;
  assign N700 = N698 & N699;
  assign N701 = N700 & N810;
  assign N702 = N701 & N259;
  assign N703 = N270 & last_r[2];
  assign N704 = N272 & N273;
  assign N705 = N258 & N259;
  assign N706 = N703 & N704;
  assign N707 = N706 & N916;
  assign N708 = N707 & N705;
  assign N709 = N270 & last_r[2];
  assign N710 = N272 & N273;
  assign N711 = N709 & N710;
  assign N712 = N819 & N259;
  assign N713 = N711 & N1027;
  assign N714 = N713 & N712;
  assign N715 = N270 & last_r[2];
  assign N716 = N272 & N273;
  assign N717 = N715 & N716;
  assign N718 = N926 & N705;
  assign N719 = N717 & N1127;
  assign N720 = N719 & N718;
  assign N721 = N270 & last_r[2];
  assign N722 = N272 & N273;
  assign N723 = N721 & N722;
  assign N724 = N723 & N1242;
  assign N725 = N832 & N259;
  assign N726 = N724 & N725;
  assign N727 = N270 & last_r[2];
  assign N728 = N272 & N273;
  assign N729 = N727 & N728;
  assign N730 = N729 & N1349;
  assign N731 = N939 & N705;
  assign N732 = N730 & N731;
  assign N733 = last_r[3] | N271;
  assign N734 = last_r[1] | last_r[0];
  assign N735 = N733 | N734;
  assign N736 = N843 | reqs_i[5];
  assign N737 = N735 | N643;
  assign N738 = N1051 | N736;
  assign N739 = N737 | N738;
  assign N742 = N270 & last_r[2];
  assign N743 = N272 & N273;
  assign N744 = N741 & N1564;
  assign N745 = N1552 & N1451;
  assign N746 = N259 & reqs_i[0];
  assign N747 = N742 & N743;
  assign N748 = N744 & N745;
  assign N749 = N1150 & N1037;
  assign N750 = N819 & N746;
  assign N751 = N747 & N748;
  assign N752 = N749 & N750;
  assign N753 = N751 & N752;
  assign N754 = N270 & last_r[2];
  assign N755 = N272 & N273;
  assign N756 = N259 & reqs_i[1];
  assign N757 = N754 & N755;
  assign N758 = N819 & N756;
  assign N759 = N757 & N748;
  assign N760 = N749 & N758;
  assign N761 = N759 & N760;
  assign N762 = N761 & N560;
  assign N763 = N270 & last_r[2];
  assign N764 = N272 & N273;
  assign N765 = N259 & reqs_i[2];
  assign N766 = N278 & N560;
  assign N767 = N763 & N764;
  assign N768 = N819 & N765;
  assign N769 = N767 & N748;
  assign N770 = N749 & N768;
  assign N771 = N769 & N770;
  assign N772 = N771 & N766;
  assign N773 = N270 & last_r[2];
  assign N774 = N272 & N273;
  assign N775 = N259 & reqs_i[3];
  assign N776 = N773 & N774;
  assign N777 = N819 & N775;
  assign N778 = N359 & N560;
  assign N779 = N776 & N748;
  assign N780 = N749 & N777;
  assign N781 = N779 & N780;
  assign N782 = N781 & N778;
  assign N783 = last_r[3] | N271;
  assign N784 = last_r[1] | last_r[0];
  assign N785 = reqs_i[5] | N260;
  assign N786 = N783 | N784;
  assign N787 = N843 | N785;
  assign N788 = N786 | N377;
  assign N789 = N1051 | N787;
  assign N790 = N788 | N789;
  assign N791 = N790 | N1953;
  assign N793 = N270 & last_r[2];
  assign N794 = N272 & last_r[0];
  assign N795 = N793 & N794;
  assign N796 = N795 & reqs_i[6];
  assign N797 = N270 & last_r[2];
  assign N798 = N272 & last_r[0];
  assign N799 = reqs_i[7] & N258;
  assign N800 = N797 & N798;
  assign N801 = N800 & N799;
  assign N802 = N270 & last_r[2];
  assign N803 = N272 & last_r[0];
  assign N804 = N802 & N803;
  assign N805 = N905 & N258;
  assign N806 = N804 & N805;
  assign N807 = N270 & last_r[2];
  assign N808 = N272 & last_r[0];
  assign N809 = N807 & N808;
  assign N810 = N1016 & N819;
  assign N811 = N809 & N810;
  assign N812 = N270 & last_r[2];
  assign N813 = N272 & last_r[0];
  assign N814 = N812 & N813;
  assign N815 = N814 & N916;
  assign N816 = N815 & N258;
  assign N817 = N270 & last_r[2];
  assign N818 = N272 & last_r[0];
  assign N819 = N918 & N258;
  assign N820 = N817 & N818;
  assign N821 = N820 & N1027;
  assign N822 = N821 & N819;
  assign N823 = N270 & last_r[2];
  assign N824 = N272 & last_r[0];
  assign N825 = N823 & N824;
  assign N826 = N926 & N258;
  assign N827 = N825 & N1127;
  assign N828 = N827 & N826;
  assign N829 = N270 & last_r[2];
  assign N830 = N272 & last_r[0];
  assign N831 = N829 & N830;
  assign N832 = N1037 & N819;
  assign N833 = N831 & N1242;
  assign N834 = N833 & N832;
  assign N835 = N270 & last_r[2];
  assign N836 = N272 & last_r[0];
  assign N837 = N835 & N836;
  assign N838 = N837 & N1349;
  assign N839 = N939 & N258;
  assign N840 = N838 & N839;
  assign N841 = last_r[3] | N271;
  assign N842 = last_r[1] | N273;
  assign N843 = reqs_i[7] | reqs_i[6];
  assign N844 = N841 | N842;
  assign N845 = N844 | N643;
  assign N846 = N1051 | N843;
  assign N847 = N845 | N846;
  assign N849 = N270 & last_r[2];
  assign N850 = N272 & last_r[0];
  assign N851 = N849 & N850;
  assign N852 = N819 & reqs_i[0];
  assign N853 = N851 & N748;
  assign N854 = N749 & N852;
  assign N855 = N853 & N854;
  assign N856 = N270 & last_r[2];
  assign N857 = N272 & last_r[0];
  assign N858 = N856 & N857;
  assign N859 = N819 & N1476;
  assign N860 = N858 & N748;
  assign N861 = N749 & N859;
  assign N862 = N860 & N861;
  assign N863 = N270 & last_r[2];
  assign N864 = N272 & last_r[0];
  assign N865 = N863 & N864;
  assign N866 = N819 & N664;
  assign N867 = N865 & N748;
  assign N868 = N749 & N866;
  assign N869 = N867 & N868;
  assign N870 = N869 & N560;
  assign N871 = N270 & last_r[2];
  assign N872 = N272 & last_r[0];
  assign N873 = N278 & N560;
  assign N874 = N871 & N872;
  assign N875 = N819 & N389;
  assign N876 = N874 & N748;
  assign N877 = N749 & N875;
  assign N878 = N876 & N877;
  assign N879 = N878 & N873;
  assign N880 = N270 & last_r[2];
  assign N881 = N272 & last_r[0];
  assign N882 = N880 & N881;
  assign N883 = N819 & N486;
  assign N884 = N359 & N560;
  assign N885 = N882 & N748;
  assign N886 = N749 & N883;
  assign N887 = N885 & N886;
  assign N888 = N887 & N884;
  assign N889 = last_r[3] | N271;
  assign N890 = last_r[1] | N273;
  assign N891 = N259 | reqs_i[4];
  assign N892 = N889 | N890;
  assign N893 = N843 | N891;
  assign N894 = N892 | N377;
  assign N895 = N1051 | N893;
  assign N896 = N894 | N895;
  assign N897 = N896 | N1953;
  assign N899 = N270 & last_r[2];
  assign N900 = last_r[1] & N273;
  assign N901 = N899 & N900;
  assign N902 = N901 & reqs_i[7];
  assign N903 = N270 & last_r[2];
  assign N904 = last_r[1] & N273;
  assign N905 = reqs_i[8] & N918;
  assign N906 = N903 & N904;
  assign N907 = N906 & N905;
  assign N908 = N270 & last_r[2];
  assign N909 = last_r[1] & N273;
  assign N910 = N908 & N909;
  assign N911 = N1016 & N918;
  assign N912 = N910 & N911;
  assign N913 = N270 & last_r[2];
  assign N914 = last_r[1] & N273;
  assign N915 = N913 & N914;
  assign N916 = N1116 & N926;
  assign N917 = N915 & N916;
  assign N919 = N270 & last_r[2];
  assign N920 = last_r[1] & N273;
  assign N921 = N919 & N920;
  assign N922 = N921 & N1027;
  assign N923 = N922 & N918;
  assign N924 = N270 & last_r[2];
  assign N925 = last_r[1] & N273;
  assign N926 = N1029 & N918;
  assign N927 = N924 & N925;
  assign N928 = N927 & N1127;
  assign N929 = N928 & N926;
  assign N930 = N270 & last_r[2];
  assign N931 = last_r[1] & N273;
  assign N932 = N930 & N931;
  assign N933 = N1037 & N918;
  assign N934 = N932 & N1242;
  assign N935 = N934 & N933;
  assign N936 = N270 & last_r[2];
  assign N937 = last_r[1] & N273;
  assign N938 = N936 & N937;
  assign N939 = N1137 & N926;
  assign N940 = N938 & N1349;
  assign N941 = N940 & N939;
  assign N942 = last_r[3] | N271;
  assign N943 = N272 | last_r[0];
  assign N944 = N942 | N943;
  assign N945 = N944 | N1466;
  assign N946 = N1051 | reqs_i[7];
  assign N947 = N945 | N946;
  assign N949 = N270 & last_r[2];
  assign N950 = last_r[1] & N273;
  assign N951 = N918 & reqs_i[0];
  assign N952 = N949 & N950;
  assign N953 = N1567 & N745;
  assign N954 = N952 & N953;
  assign N955 = N749 & N951;
  assign N956 = N954 & N955;
  assign N957 = N270 & last_r[2];
  assign N958 = last_r[1] & N273;
  assign N959 = N918 & reqs_i[1];
  assign N960 = N957 & N958;
  assign N961 = N959 & N560;
  assign N962 = N960 & N953;
  assign N963 = N749 & N961;
  assign N964 = N962 & N963;
  assign N965 = N270 & last_r[2];
  assign N966 = last_r[1] & N273;
  assign N967 = N918 & reqs_i[2];
  assign N968 = N965 & N966;
  assign N969 = N967 & N873;
  assign N970 = N968 & N953;
  assign N971 = N749 & N969;
  assign N972 = N970 & N971;
  assign N973 = N270 & last_r[2];
  assign N974 = last_r[1] & N273;
  assign N975 = N918 & reqs_i[3];
  assign N976 = N973 & N974;
  assign N977 = N975 & N359;
  assign N978 = N976 & N953;
  assign N979 = N749 & N977;
  assign N980 = N978 & N979;
  assign N981 = N980 & N560;
  assign N982 = N270 & last_r[2];
  assign N983 = last_r[1] & N273;
  assign N984 = N918 & reqs_i[4];
  assign N985 = N982 & N983;
  assign N986 = N984 & N409;
  assign N987 = N985 & N953;
  assign N988 = N749 & N986;
  assign N989 = N987 & N988;
  assign N990 = N989 & N873;
  assign N991 = N270 & last_r[2];
  assign N992 = last_r[1] & N273;
  assign N993 = N918 & reqs_i[5];
  assign N994 = N991 & N992;
  assign N995 = N993 & N506;
  assign N996 = N994 & N953;
  assign N997 = N749 & N995;
  assign N998 = N996 & N997;
  assign N999 = N998 & N884;
  assign N1000 = last_r[3] | N271;
  assign N1001 = N272 | last_r[0];
  assign N1002 = reqs_i[7] | N258;
  assign N1003 = N1000 | N1001;
  assign N1004 = N1002 | N641;
  assign N1005 = N1003 | N377;
  assign N1006 = N1051 | N1004;
  assign N1007 = N1005 | N1006;
  assign N1008 = N1007 | N1953;
  assign N1010 = N270 & last_r[2];
  assign N1011 = last_r[1] & last_r[0];
  assign N1012 = N1010 & N1011;
  assign N1013 = N1012 & reqs_i[8];
  assign N1014 = N270 & last_r[2];
  assign N1015 = last_r[1] & last_r[0];
  assign N1016 = reqs_i[9] & N1029;
  assign N1017 = N1014 & N1015;
  assign N1018 = N1017 & N1016;
  assign N1019 = N270 & last_r[2];
  assign N1020 = last_r[1] & last_r[0];
  assign N1021 = N1019 & N1020;
  assign N1022 = N1116 & N1029;
  assign N1023 = N1021 & N1022;
  assign N1024 = N270 & last_r[2];
  assign N1025 = last_r[1] & last_r[0];
  assign N1026 = N1024 & N1025;
  assign N1027 = N1231 & N1037;
  assign N1028 = N1026 & N1027;
  assign N1030 = N270 & last_r[2];
  assign N1031 = last_r[1] & last_r[0];
  assign N1032 = N1030 & N1031;
  assign N1033 = N1032 & N1127;
  assign N1034 = N1033 & N1029;
  assign N1035 = N270 & last_r[2];
  assign N1036 = last_r[1] & last_r[0];
  assign N1037 = N1129 & N1029;
  assign N1038 = N1035 & N1036;
  assign N1039 = N1038 & N1242;
  assign N1040 = N1039 & N1037;
  assign N1041 = N270 & last_r[2];
  assign N1042 = last_r[1] & last_r[0];
  assign N1043 = N1041 & N1042;
  assign N1044 = N1137 & N1029;
  assign N1045 = N1043 & N1349;
  assign N1046 = N1045 & N1044;
  assign N1047 = last_r[3] | N271;
  assign N1048 = N272 | N273;
  assign N1049 = reqs_i[9] | reqs_i[8];
  assign N1050 = N1047 | N1048;
  assign N1051 = N1252 | N1049;
  assign N1052 = N1050 | N1466;
  assign N1053 = N1052 | N1051;
  assign N1055 = N270 & last_r[2];
  assign N1056 = last_r[1] & last_r[0];
  assign N1057 = N1055 & N1056;
  assign N1058 = N1057 & N953;
  assign N1059 = N749 & reqs_i[0];
  assign N1060 = N1058 & N1059;
  assign N1061 = N270 & last_r[2];
  assign N1062 = last_r[1] & last_r[0];
  assign N1063 = N1061 & N1062;
  assign N1064 = N1063 & N953;
  assign N1065 = N749 & N1476;
  assign N1066 = N1064 & N1065;
  assign N1067 = N270 & last_r[2];
  assign N1068 = last_r[1] & last_r[0];
  assign N1069 = N1067 & N1068;
  assign N1070 = N1069 & N953;
  assign N1071 = N749 & N1483;
  assign N1072 = N1070 & N1071;
  assign N1073 = N270 & last_r[2];
  assign N1074 = last_r[1] & last_r[0];
  assign N1075 = N1073 & N1074;
  assign N1076 = N1075 & N953;
  assign N1077 = N749 & N1489;
  assign N1078 = N1076 & N1077;
  assign N1079 = N270 & last_r[2];
  assign N1080 = last_r[1] & last_r[0];
  assign N1081 = N1079 & N1080;
  assign N1082 = N1081 & N953;
  assign N1083 = N749 & N1495;
  assign N1084 = N1082 & N1083;
  assign N1085 = N1084 & N560;
  assign N1086 = N270 & last_r[2];
  assign N1087 = last_r[1] & last_r[0];
  assign N1088 = N1086 & N1087;
  assign N1089 = N1088 & N953;
  assign N1090 = N749 & N400;
  assign N1091 = N1089 & N1090;
  assign N1092 = N1091 & N873;
  assign N1093 = N270 & last_r[2];
  assign N1094 = last_r[1] & last_r[0];
  assign N1095 = N1093 & N1094;
  assign N1096 = N1095 & N953;
  assign N1097 = N749 & N497;
  assign N1098 = N1096 & N1097;
  assign N1099 = N1098 & N884;
  assign N1100 = last_r[3] | N271;
  assign N1101 = N272 | N273;
  assign N1102 = N918 | reqs_i[6];
  assign N1103 = N1100 | N1101;
  assign N1104 = N1102 | N641;
  assign N1105 = N1103 | N377;
  assign N1106 = N1051 | N1104;
  assign N1107 = N1105 | N1106;
  assign N1108 = N1107 | N1953;
  assign N1110 = last_r[3] & N271;
  assign N1111 = N272 & N273;
  assign N1112 = N1110 & N1111;
  assign N1113 = N1112 & reqs_i[9];
  assign N1114 = last_r[3] & N271;
  assign N1115 = N272 & N273;
  assign N1116 = reqs_i[10] & N1129;
  assign N1117 = N1114 & N1115;
  assign N1118 = N1117 & N1116;
  assign N1119 = last_r[3] & N271;
  assign N1120 = N272 & N273;
  assign N1121 = N1119 & N1120;
  assign N1122 = N1231 & N1129;
  assign N1123 = N1121 & N1122;
  assign N1124 = last_r[3] & N271;
  assign N1125 = N272 & N273;
  assign N1126 = N1124 & N1125;
  assign N1127 = N1337 & N1137;
  assign N1128 = N1126 & N1127;
  assign N1130 = last_r[3] & N271;
  assign N1131 = N272 & N273;
  assign N1132 = N1130 & N1131;
  assign N1133 = N1132 & N1242;
  assign N1134 = N1133 & N1129;
  assign N1135 = last_r[3] & N271;
  assign N1136 = N272 & N273;
  assign N1137 = N1244 & N1129;
  assign N1138 = N1135 & N1136;
  assign N1139 = N1138 & N1349;
  assign N1140 = N1139 & N1137;
  assign N1141 = N270 | last_r[2];
  assign N1142 = last_r[1] | last_r[0];
  assign N1143 = N1141 | N1142;
  assign N1144 = N1252 | reqs_i[9];
  assign N1145 = N1143 | N1466;
  assign N1146 = N1145 | N1144;
  assign N1148 = last_r[3] & N271;
  assign N1149 = N272 & N273;
  assign N1150 = N1357 & N1244;
  assign N1151 = N1129 & reqs_i[0];
  assign N1152 = N1148 & N1149;
  assign N1153 = N1150 & N1151;
  assign N1154 = N1152 & N953;
  assign N1155 = N1154 & N1153;
  assign N1156 = last_r[3] & N271;
  assign N1157 = N272 & N273;
  assign N1158 = N1129 & reqs_i[1];
  assign N1159 = N1156 & N1157;
  assign N1160 = N1150 & N1158;
  assign N1161 = N1159 & N953;
  assign N1162 = N1160 & N560;
  assign N1163 = N1161 & N1162;
  assign N1164 = last_r[3] & N271;
  assign N1165 = N272 & N273;
  assign N1166 = N1129 & reqs_i[2];
  assign N1167 = N1164 & N1165;
  assign N1168 = N1150 & N1166;
  assign N1169 = N1167 & N953;
  assign N1170 = N1168 & N873;
  assign N1171 = N1169 & N1170;
  assign N1172 = last_r[3] & N271;
  assign N1173 = N272 & N273;
  assign N1174 = N1129 & reqs_i[3];
  assign N1175 = N1172 & N1173;
  assign N1176 = N1150 & N1174;
  assign N1177 = N1175 & N953;
  assign N1178 = N1176 & N884;
  assign N1179 = N1177 & N1178;
  assign N1180 = last_r[3] & N271;
  assign N1181 = N272 & N273;
  assign N1182 = N1129 & reqs_i[4];
  assign N1183 = N1180 & N1181;
  assign N1184 = N1150 & N1182;
  assign N1185 = N1183 & N953;
  assign N1186 = N1184 & N1598;
  assign N1187 = N1185 & N1186;
  assign N1188 = last_r[3] & N271;
  assign N1189 = N272 & N273;
  assign N1190 = N1129 & reqs_i[5];
  assign N1191 = N1188 & N1189;
  assign N1192 = N1150 & N1190;
  assign N1193 = N1191 & N953;
  assign N1194 = N1192 & N323;
  assign N1195 = N1193 & N1194;
  assign N1196 = N1195 & N560;
  assign N1197 = last_r[3] & N271;
  assign N1198 = N272 & N273;
  assign N1199 = N1129 & reqs_i[6];
  assign N1200 = N1197 & N1198;
  assign N1201 = N1150 & N1199;
  assign N1202 = N1200 & N953;
  assign N1203 = N1201 & N422;
  assign N1204 = N1202 & N1203;
  assign N1205 = N1204 & N873;
  assign N1206 = last_r[3] & N271;
  assign N1207 = N272 & N273;
  assign N1208 = N1129 & reqs_i[7];
  assign N1209 = N1206 & N1207;
  assign N1210 = N1150 & N1208;
  assign N1211 = N1209 & N953;
  assign N1212 = N1210 & N519;
  assign N1213 = N1211 & N1212;
  assign N1214 = N1213 & N884;
  assign N1215 = N270 | last_r[2];
  assign N1216 = last_r[1] | last_r[0];
  assign N1217 = reqs_i[9] | N1029;
  assign N1218 = N1215 | N1216;
  assign N1219 = N1252 | N1217;
  assign N1220 = N1218 | N377;
  assign N1221 = N1219 | N644;
  assign N1222 = N1220 | N1221;
  assign N1223 = N1222 | N1953;
  assign N1225 = last_r[3] & N271;
  assign N1226 = N272 & last_r[0];
  assign N1227 = N1225 & N1226;
  assign N1228 = N1227 & reqs_i[10];
  assign N1229 = last_r[3] & N271;
  assign N1230 = N272 & last_r[0];
  assign N1231 = reqs_i[11] & N1244;
  assign N1232 = N1229 & N1230;
  assign N1233 = N1232 & N1231;
  assign N1234 = last_r[3] & N271;
  assign N1235 = N272 & last_r[0];
  assign N1236 = N1234 & N1235;
  assign N1237 = N1337 & N1244;
  assign N1238 = N1236 & N1237;
  assign N1239 = last_r[3] & N271;
  assign N1240 = N272 & last_r[0];
  assign N1241 = N1239 & N1240;
  assign N1242 = N1454 & N1150;
  assign N1243 = N1241 & N1242;
  assign N1245 = last_r[3] & N271;
  assign N1246 = N272 & last_r[0];
  assign N1247 = N1245 & N1246;
  assign N1248 = N1247 & N1349;
  assign N1249 = N1248 & N1244;
  assign N1250 = N270 | last_r[2];
  assign N1251 = last_r[1] | N273;
  assign N1252 = reqs_i[11] | reqs_i[10];
  assign N1253 = N1250 | N1251;
  assign N1254 = N1253 | N1466;
  assign N1255 = N1254 | N1252;
  assign N1257 = last_r[3] & N271;
  assign N1258 = N272 & last_r[0];
  assign N1259 = N1257 & N1258;
  assign N1260 = N1150 & reqs_i[0];
  assign N1261 = N1259 & N953;
  assign N1262 = N1261 & N1260;
  assign N1263 = last_r[3] & N271;
  assign N1264 = N272 & last_r[0];
  assign N1265 = N1263 & N1264;
  assign N1266 = N1150 & N1476;
  assign N1267 = N1265 & N953;
  assign N1268 = N1267 & N1266;
  assign N1269 = last_r[3] & N271;
  assign N1270 = N272 & last_r[0];
  assign N1271 = N1269 & N1270;
  assign N1272 = N1150 & N664;
  assign N1273 = N1271 & N953;
  assign N1274 = N1272 & N560;
  assign N1275 = N1273 & N1274;
  assign N1276 = last_r[3] & N271;
  assign N1277 = N272 & last_r[0];
  assign N1278 = N1276 & N1277;
  assign N1279 = N1150 & N389;
  assign N1280 = N1278 & N953;
  assign N1281 = N1279 & N873;
  assign N1282 = N1280 & N1281;
  assign N1283 = last_r[3] & N271;
  assign N1284 = N272 & last_r[0];
  assign N1285 = N1283 & N1284;
  assign N1286 = N1150 & N486;
  assign N1287 = N1285 & N953;
  assign N1288 = N1286 & N884;
  assign N1289 = N1287 & N1288;
  assign N1290 = last_r[3] & N271;
  assign N1291 = N272 & last_r[0];
  assign N1292 = N1290 & N1291;
  assign N1293 = N1150 & N584;
  assign N1294 = N1292 & N953;
  assign N1295 = N1293 & N1598;
  assign N1296 = N1294 & N1295;
  assign N1297 = last_r[3] & N271;
  assign N1298 = N272 & last_r[0];
  assign N1299 = N1297 & N1298;
  assign N1300 = N1150 & N685;
  assign N1301 = N1299 & N953;
  assign N1302 = N1300 & N323;
  assign N1303 = N1301 & N1302;
  assign N1304 = N1303 & N560;
  assign N1305 = last_r[3] & N271;
  assign N1306 = N272 & last_r[0];
  assign N1307 = N1305 & N1306;
  assign N1308 = N1150 & N799;
  assign N1309 = N1307 & N953;
  assign N1310 = N1308 & N422;
  assign N1311 = N1309 & N1310;
  assign N1312 = N1311 & N873;
  assign N1313 = last_r[3] & N271;
  assign N1314 = N272 & last_r[0];
  assign N1315 = N1313 & N1314;
  assign N1316 = N1150 & N905;
  assign N1317 = N1315 & N953;
  assign N1318 = N1316 & N519;
  assign N1319 = N1317 & N1318;
  assign N1320 = N1319 & N884;
  assign N1321 = N270 | last_r[2];
  assign N1322 = last_r[1] | N273;
  assign N1323 = N1129 | reqs_i[8];
  assign N1324 = N1321 | N1322;
  assign N1325 = N1252 | N1323;
  assign N1326 = N1324 | N377;
  assign N1327 = N1325 | N644;
  assign N1328 = N1326 | N1327;
  assign N1329 = N1328 | N1953;
  assign N1331 = last_r[3] & N271;
  assign N1332 = last_r[1] & N273;
  assign N1333 = N1331 & N1332;
  assign N1334 = N1333 & reqs_i[11];
  assign N1335 = last_r[3] & N271;
  assign N1336 = last_r[1] & N273;
  assign N1337 = reqs_i[12] & N1357;
  assign N1338 = N1335 & N1336;
  assign N1339 = N1338 & N1337;
  assign N1340 = last_r[3] & N271;
  assign N1341 = last_r[1] & N273;
  assign N1342 = N1340 & N1341;
  assign N1343 = N1454 & N1357;
  assign N1344 = N1342 & N1343;
  assign N1345 = last_r[3] & N271;
  assign N1346 = last_r[1] & N273;
  assign N1347 = N1451 & N1357;
  assign N1348 = N1345 & N1346;
  assign N1349 = N1555 & N1347;
  assign N1350 = N1348 & N1349;
  assign N1351 = N270 | last_r[2];
  assign N1352 = N272 | last_r[0];
  assign N1353 = N1351 | N1352;
  assign N1354 = N1353 | N1466;
  assign N1355 = N1354 | reqs_i[11];
  assign N1358 = last_r[3] & N271;
  assign N1359 = last_r[1] & N273;
  assign N1360 = N1357 & reqs_i[0];
  assign N1361 = N1358 & N1359;
  assign N1362 = N1361 & N953;
  assign N1363 = N1362 & N1360;
  assign N1364 = last_r[3] & N271;
  assign N1365 = last_r[1] & N273;
  assign N1366 = N1357 & reqs_i[1];
  assign N1367 = N1364 & N1365;
  assign N1368 = N1366 & N560;
  assign N1369 = N1367 & N953;
  assign N1370 = N1369 & N1368;
  assign N1371 = last_r[3] & N271;
  assign N1372 = last_r[1] & N273;
  assign N1373 = N1357 & reqs_i[2];
  assign N1374 = N1371 & N1372;
  assign N1375 = N1373 & N873;
  assign N1376 = N1374 & N953;
  assign N1377 = N1376 & N1375;
  assign N1378 = last_r[3] & N271;
  assign N1379 = last_r[1] & N273;
  assign N1380 = N1357 & reqs_i[3];
  assign N1381 = N1378 & N1379;
  assign N1382 = N1380 & N359;
  assign N1383 = N1381 & N953;
  assign N1384 = N1382 & N560;
  assign N1385 = N1383 & N1384;
  assign N1386 = last_r[3] & N271;
  assign N1387 = last_r[1] & N273;
  assign N1388 = N1357 & reqs_i[4];
  assign N1389 = N1386 & N1387;
  assign N1390 = N1388 & N409;
  assign N1391 = N1389 & N953;
  assign N1392 = N1390 & N873;
  assign N1393 = N1391 & N1392;
  assign N1394 = last_r[3] & N271;
  assign N1395 = last_r[1] & N273;
  assign N1396 = N1357 & reqs_i[5];
  assign N1397 = N1394 & N1395;
  assign N1398 = N1396 & N506;
  assign N1399 = N1397 & N953;
  assign N1400 = N1398 & N884;
  assign N1401 = N1399 & N1400;
  assign N1402 = last_r[3] & N271;
  assign N1403 = last_r[1] & N273;
  assign N1404 = N1357 & reqs_i[6];
  assign N1405 = N1402 & N1403;
  assign N1406 = N1404 & N604;
  assign N1407 = N1405 & N953;
  assign N1408 = N1406 & N1598;
  assign N1409 = N1407 & N1408;
  assign N1410 = last_r[3] & N271;
  assign N1411 = last_r[1] & N273;
  assign N1412 = N1357 & reqs_i[7];
  assign N1413 = N1410 & N1411;
  assign N1414 = N1412 & N705;
  assign N1415 = N1413 & N953;
  assign N1416 = N1414 & N323;
  assign N1417 = N1415 & N1416;
  assign N1418 = N1417 & N560;
  assign N1419 = last_r[3] & N271;
  assign N1420 = last_r[1] & N273;
  assign N1421 = N1357 & reqs_i[8];
  assign N1422 = N1419 & N1420;
  assign N1423 = N1421 & N819;
  assign N1424 = N1422 & N953;
  assign N1425 = N1423 & N422;
  assign N1426 = N1424 & N1425;
  assign N1427 = N1426 & N873;
  assign N1428 = last_r[3] & N271;
  assign N1429 = last_r[1] & N273;
  assign N1430 = N1357 & reqs_i[9];
  assign N1431 = N1428 & N1429;
  assign N1432 = N1430 & N926;
  assign N1433 = N1431 & N953;
  assign N1434 = N1432 & N519;
  assign N1435 = N1433 & N1434;
  assign N1436 = N1435 & N884;
  assign N1437 = N270 | last_r[2];
  assign N1438 = N272 | last_r[0];
  assign N1439 = reqs_i[11] | N1244;
  assign N1440 = N1437 | N1438;
  assign N1441 = N1439 | N1049;
  assign N1442 = N1440 | N377;
  assign N1443 = N1441 | N644;
  assign N1444 = N1442 | N1443;
  assign N1445 = N1444 | N1953;
  assign N1447 = last_r[3] & N271;
  assign N1448 = last_r[1] & last_r[0];
  assign N1449 = N1447 & N1448;
  assign N1450 = N1449 & reqs_i[12];
  assign N1452 = last_r[3] & N271;
  assign N1453 = last_r[1] & last_r[0];
  assign N1454 = reqs_i[13] & N1451;
  assign N1455 = N1452 & N1453;
  assign N1456 = N1455 & N1454;
  assign N1457 = last_r[3] & N271;
  assign N1458 = last_r[1] & last_r[0];
  assign N1459 = N1457 & N1458;
  assign N1460 = N1555 & N1451;
  assign N1461 = N1459 & N1460;
  assign N1462 = N270 | last_r[2];
  assign N1463 = N272 | N273;
  assign N1464 = reqs_i[13] | reqs_i[12];
  assign N1465 = N1462 | N1463;
  assign N1466 = N1672 | N1464;
  assign N1467 = N1465 | N1466;
  assign N1469 = last_r[3] & N271;
  assign N1470 = last_r[1] & last_r[0];
  assign N1471 = N1469 & N1470;
  assign N1472 = N1471 & N953;
  assign N1473 = N1472 & reqs_i[0];
  assign N1474 = last_r[3] & N271;
  assign N1475 = last_r[1] & last_r[0];
  assign N1476 = reqs_i[1] & N560;
  assign N1477 = N1474 & N1475;
  assign N1478 = N1477 & N953;
  assign N1479 = N1478 & N1476;
  assign N1480 = last_r[3] & N271;
  assign N1481 = last_r[1] & last_r[0];
  assign N1482 = N1480 & N1481;
  assign N1483 = N664 & N560;
  assign N1484 = N1482 & N953;
  assign N1485 = N1484 & N1483;
  assign N1486 = last_r[3] & N271;
  assign N1487 = last_r[1] & last_r[0];
  assign N1488 = N1486 & N1487;
  assign N1489 = N389 & N873;
  assign N1490 = N1488 & N953;
  assign N1491 = N1490 & N1489;
  assign N1492 = last_r[3] & N271;
  assign N1493 = last_r[1] & last_r[0];
  assign N1494 = N1492 & N1493;
  assign N1495 = N486 & N359;
  assign N1496 = N1494 & N953;
  assign N1497 = N1495 & N560;
  assign N1498 = N1496 & N1497;
  assign N1499 = last_r[3] & N271;
  assign N1500 = last_r[1] & last_r[0];
  assign N1501 = N1499 & N1500;
  assign N1502 = N1501 & N953;
  assign N1503 = N400 & N873;
  assign N1504 = N1502 & N1503;
  assign N1505 = last_r[3] & N271;
  assign N1506 = last_r[1] & last_r[0];
  assign N1507 = N1505 & N1506;
  assign N1508 = N1507 & N953;
  assign N1509 = N497 & N884;
  assign N1510 = N1508 & N1509;
  assign N1511 = last_r[3] & N271;
  assign N1512 = last_r[1] & last_r[0];
  assign N1513 = N1511 & N1512;
  assign N1514 = N1513 & N953;
  assign N1515 = N595 & N1598;
  assign N1516 = N1514 & N1515;
  assign N1517 = last_r[3] & N271;
  assign N1518 = last_r[1] & last_r[0];
  assign N1519 = N1517 & N1518;
  assign N1520 = N1519 & N953;
  assign N1521 = N696 & N323;
  assign N1522 = N1520 & N1521;
  assign N1523 = N1522 & N560;
  assign N1524 = last_r[3] & N271;
  assign N1525 = last_r[1] & last_r[0];
  assign N1526 = N1524 & N1525;
  assign N1527 = N1526 & N953;
  assign N1528 = N810 & N422;
  assign N1529 = N1527 & N1528;
  assign N1530 = N1529 & N873;
  assign N1531 = last_r[3] & N271;
  assign N1532 = last_r[1] & last_r[0];
  assign N1533 = N1531 & N1532;
  assign N1534 = N1533 & N953;
  assign N1535 = N916 & N519;
  assign N1536 = N1534 & N1535;
  assign N1537 = N1536 & N884;
  assign N1538 = N270 | last_r[2];
  assign N1539 = N272 | N273;
  assign N1540 = N1357 | reqs_i[10];
  assign N1541 = N1538 | N1539;
  assign N1542 = N1540 | N1049;
  assign N1543 = N1541 | N377;
  assign N1544 = N1542 | N644;
  assign N1545 = N1543 | N1544;
  assign N1546 = N1545 | N1953;
  assign N1548 = last_r[3] & last_r[2];
  assign N1549 = N272 & N273;
  assign N1550 = N1548 & N1549;
  assign N1551 = N1550 & reqs_i[13];
  assign N1553 = last_r[3] & last_r[2];
  assign N1554 = N272 & N273;
  assign N1555 = reqs_i[14] & N1552;
  assign N1556 = N1553 & N1554;
  assign N1557 = N1556 & N1555;
  assign N1558 = N270 | N271;
  assign N1559 = last_r[1] | last_r[0];
  assign N1560 = N1558 | N1559;
  assign N1561 = N1672 | reqs_i[13];
  assign N1562 = N1560 | N1561;
  assign N1565 = last_r[3] & last_r[2];
  assign N1566 = N272 & N273;
  assign N1567 = N741 & N1564;
  assign N1568 = N1552 & reqs_i[0];
  assign N1569 = N1565 & N1566;
  assign N1570 = N1567 & N1568;
  assign N1571 = N1569 & N1570;
  assign N1572 = last_r[3] & last_r[2];
  assign N1573 = N272 & N273;
  assign N1574 = N1552 & reqs_i[1];
  assign N1575 = N1572 & N1573;
  assign N1576 = N1567 & N1574;
  assign N1577 = N1575 & N1576;
  assign N1578 = N1577 & N560;
  assign N1579 = last_r[3] & last_r[2];
  assign N1580 = N272 & N273;
  assign N1581 = N1552 & reqs_i[2];
  assign N1582 = N1579 & N1580;
  assign N1583 = N1567 & N1581;
  assign N1584 = N1582 & N1583;
  assign N1585 = N1584 & N873;
  assign N1586 = last_r[3] & last_r[2];
  assign N1587 = N272 & N273;
  assign N1588 = N1552 & reqs_i[3];
  assign N1589 = N1586 & N1587;
  assign N1590 = N1567 & N1588;
  assign N1591 = N1589 & N1590;
  assign N1592 = N1591 & N884;
  assign N1593 = last_r[3] & last_r[2];
  assign N1594 = N272 & N273;
  assign N1595 = N1552 & reqs_i[4];
  assign N1596 = N1593 & N1594;
  assign N1597 = N1567 & N1595;
  assign N1598 = N409 & N873;
  assign N1599 = N1596 & N1597;
  assign N1600 = N1599 & N1598;
  assign N1601 = last_r[3] & last_r[2];
  assign N1602 = N272 & N273;
  assign N1603 = N1552 & reqs_i[5];
  assign N1604 = N1601 & N1602;
  assign N1605 = N1567 & N1603;
  assign N1606 = N1604 & N1605;
  assign N1607 = N323 & N560;
  assign N1608 = N1606 & N1607;
  assign N1609 = last_r[3] & last_r[2];
  assign N1610 = N272 & N273;
  assign N1611 = N1552 & reqs_i[6];
  assign N1612 = N1609 & N1610;
  assign N1613 = N1567 & N1611;
  assign N1614 = N1612 & N1613;
  assign N1615 = N422 & N873;
  assign N1616 = N1614 & N1615;
  assign N1617 = last_r[3] & last_r[2];
  assign N1618 = N272 & N273;
  assign N1619 = N1552 & reqs_i[7];
  assign N1620 = N1617 & N1618;
  assign N1621 = N1567 & N1619;
  assign N1622 = N1620 & N1621;
  assign N1623 = N519 & N884;
  assign N1624 = N1622 & N1623;
  assign N1625 = last_r[3] & last_r[2];
  assign N1626 = N272 & N273;
  assign N1627 = N1552 & reqs_i[8];
  assign N1628 = N1625 & N1626;
  assign N1629 = N1567 & N1627;
  assign N1630 = N1628 & N1629;
  assign N1631 = N617 & N1598;
  assign N1632 = N1630 & N1631;
  assign N1633 = last_r[3] & last_r[2];
  assign N1634 = N272 & N273;
  assign N1635 = N1552 & reqs_i[9];
  assign N1636 = N1633 & N1634;
  assign N1637 = N1567 & N1635;
  assign N1638 = N1636 & N1637;
  assign N1639 = N1638 & N349;
  assign N1640 = N1639 & N560;
  assign N1641 = last_r[3] & last_r[2];
  assign N1642 = N272 & N273;
  assign N1643 = N1552 & reqs_i[10];
  assign N1644 = N1641 & N1642;
  assign N1645 = N1567 & N1643;
  assign N1646 = N1644 & N1645;
  assign N1647 = N1646 & N447;
  assign N1648 = N1647 & N873;
  assign N1649 = last_r[3] & last_r[2];
  assign N1650 = N272 & N273;
  assign N1651 = N1552 & reqs_i[11];
  assign N1652 = N1649 & N1650;
  assign N1653 = N1567 & N1651;
  assign N1654 = N1652 & N1653;
  assign N1655 = N1654 & N544;
  assign N1656 = N1655 & N884;
  assign N1657 = N270 | N271;
  assign N1658 = last_r[1] | last_r[0];
  assign N1659 = reqs_i[13] | N1451;
  assign N1660 = N1657 | N1658;
  assign N1661 = N374 | N1659;
  assign N1662 = N1660 | N1661;
  assign N1663 = N1662 | N646;
  assign N1664 = N1663 | N1953;
  assign N1666 = last_r[3] & last_r[2];
  assign N1667 = N272 & last_r[0];
  assign N1668 = N1666 & N1667;
  assign N1669 = N1668 & reqs_i[14];
  assign N1670 = N270 | N271;
  assign N1671 = last_r[1] | N273;
  assign N1672 = N741 | reqs_i[14];
  assign N1673 = N1670 | N1671;
  assign N1674 = N1673 | N1672;
  assign N1676 = last_r[3] & last_r[2];
  assign N1677 = N272 & last_r[0];
  assign N1678 = N1676 & N1677;
  assign N1679 = N1567 & reqs_i[0];
  assign N1680 = N1678 & N1679;
  assign N1681 = last_r[3] & last_r[2];
  assign N1682 = N272 & last_r[0];
  assign N1683 = N1681 & N1682;
  assign N1684 = N1567 & N1476;
  assign N1685 = N1683 & N1684;
  assign N1686 = last_r[3] & last_r[2];
  assign N1687 = N272 & last_r[0];
  assign N1688 = N1686 & N1687;
  assign N1689 = N1567 & N664;
  assign N1690 = N1688 & N1689;
  assign N1691 = N1690 & N560;
  assign N1692 = last_r[3] & last_r[2];
  assign N1693 = N272 & last_r[0];
  assign N1694 = N1692 & N1693;
  assign N1695 = N1567 & N389;
  assign N1696 = N1694 & N1695;
  assign N1697 = N1696 & N873;
  assign N1698 = last_r[3] & last_r[2];
  assign N1699 = N272 & last_r[0];
  assign N1700 = N1698 & N1699;
  assign N1701 = N1567 & N486;
  assign N1702 = N1700 & N1701;
  assign N1703 = N1702 & N884;
  assign N1704 = last_r[3] & last_r[2];
  assign N1705 = N272 & last_r[0];
  assign N1706 = N1704 & N1705;
  assign N1707 = N1567 & N584;
  assign N1708 = N1706 & N1707;
  assign N1709 = N1708 & N1598;
  assign N1710 = last_r[3] & last_r[2];
  assign N1711 = N272 & last_r[0];
  assign N1712 = N1710 & N1711;
  assign N1713 = N1567 & N685;
  assign N1714 = N1712 & N1713;
  assign N1715 = N1714 & N1607;
  assign N1716 = last_r[3] & last_r[2];
  assign N1717 = N272 & last_r[0];
  assign N1718 = N1716 & N1717;
  assign N1719 = N1567 & N799;
  assign N1720 = N1718 & N1719;
  assign N1721 = N1720 & N1615;
  assign N1722 = last_r[3] & last_r[2];
  assign N1723 = N272 & last_r[0];
  assign N1724 = N1722 & N1723;
  assign N1725 = N1567 & N905;
  assign N1726 = N1724 & N1725;
  assign N1727 = N1726 & N1623;
  assign N1728 = last_r[3] & last_r[2];
  assign N1729 = N272 & last_r[0];
  assign N1730 = N1728 & N1729;
  assign N1731 = N1567 & N1016;
  assign N1732 = N1730 & N1731;
  assign N1733 = N1732 & N1631;
  assign N1734 = last_r[3] & last_r[2];
  assign N1735 = N272 & last_r[0];
  assign N1736 = N1734 & N1735;
  assign N1737 = N1567 & N1116;
  assign N1738 = N1736 & N1737;
  assign N1739 = N1738 & N349;
  assign N1740 = N1739 & N560;
  assign N1741 = last_r[3] & last_r[2];
  assign N1742 = N272 & last_r[0];
  assign N1743 = N1741 & N1742;
  assign N1744 = N1567 & N1231;
  assign N1745 = N1743 & N1744;
  assign N1746 = N1745 & N447;
  assign N1747 = N1746 & N873;
  assign N1748 = last_r[3] & last_r[2];
  assign N1749 = N272 & last_r[0];
  assign N1750 = N1748 & N1749;
  assign N1751 = N1567 & N1337;
  assign N1752 = N1750 & N1751;
  assign N1753 = N1752 & N544;
  assign N1754 = N1753 & N884;
  assign N1755 = N270 | N271;
  assign N1756 = last_r[1] | N273;
  assign N1757 = N1552 | reqs_i[12];
  assign N1758 = N1755 | N1756;
  assign N1759 = N374 | N1757;
  assign N1760 = N1758 | N1759;
  assign N1761 = N1760 | N646;
  assign N1762 = N1761 | N1953;
  assign N1764 = N270 | N271;
  assign N1765 = N272 | last_r[0];
  assign N1766 = N1764 | N1765;
  assign N1767 = N1766 | N741;
  assign N1769 = last_r[3] & last_r[2];
  assign N1770 = last_r[1] & N273;
  assign N1771 = N741 & reqs_i[0];
  assign N1772 = N1769 & N1770;
  assign N1773 = N1772 & N1771;
  assign N1774 = last_r[3] & last_r[2];
  assign N1775 = last_r[1] & N273;
  assign N1776 = N741 & reqs_i[1];
  assign N1777 = N1774 & N1775;
  assign N1778 = N1776 & N560;
  assign N1779 = N1777 & N1778;
  assign N1780 = last_r[3] & last_r[2];
  assign N1781 = last_r[1] & N273;
  assign N1782 = N741 & reqs_i[2];
  assign N1783 = N1780 & N1781;
  assign N1784 = N1782 & N873;
  assign N1785 = N1783 & N1784;
  assign N1786 = last_r[3] & last_r[2];
  assign N1787 = last_r[1] & N273;
  assign N1788 = N741 & reqs_i[3];
  assign N1789 = N1786 & N1787;
  assign N1790 = N1788 & N359;
  assign N1791 = N1789 & N1790;
  assign N1792 = N1791 & N560;
  assign N1793 = last_r[3] & last_r[2];
  assign N1794 = last_r[1] & N273;
  assign N1795 = N741 & reqs_i[4];
  assign N1796 = N1793 & N1794;
  assign N1797 = N1795 & N409;
  assign N1798 = N1796 & N1797;
  assign N1799 = N1798 & N873;
  assign N1800 = last_r[3] & last_r[2];
  assign N1801 = last_r[1] & N273;
  assign N1802 = N741 & reqs_i[5];
  assign N1803 = N1800 & N1801;
  assign N1804 = N1802 & N506;
  assign N1805 = N1803 & N1804;
  assign N1806 = N1805 & N884;
  assign N1807 = last_r[3] & last_r[2];
  assign N1808 = last_r[1] & N273;
  assign N1809 = N741 & reqs_i[6];
  assign N1810 = N1807 & N1808;
  assign N1811 = N1809 & N604;
  assign N1812 = N1810 & N1811;
  assign N1813 = N1812 & N1598;
  assign N1814 = last_r[3] & last_r[2];
  assign N1815 = last_r[1] & N273;
  assign N1816 = N741 & reqs_i[7];
  assign N1817 = N1814 & N1815;
  assign N1818 = N1816 & N705;
  assign N1819 = N1817 & N1818;
  assign N1820 = N1819 & N1607;
  assign N1821 = last_r[3] & last_r[2];
  assign N1822 = last_r[1] & N273;
  assign N1823 = N741 & reqs_i[8];
  assign N1824 = N1821 & N1822;
  assign N1825 = N1823 & N819;
  assign N1826 = N1824 & N1825;
  assign N1827 = N1826 & N1615;
  assign N1828 = last_r[3] & last_r[2];
  assign N1829 = last_r[1] & N273;
  assign N1830 = N741 & reqs_i[9];
  assign N1831 = N1828 & N1829;
  assign N1832 = N1830 & N926;
  assign N1833 = N1831 & N1832;
  assign N1834 = N1833 & N1623;
  assign N1835 = last_r[3] & last_r[2];
  assign N1836 = last_r[1] & N273;
  assign N1837 = N741 & reqs_i[10];
  assign N1838 = N1835 & N1836;
  assign N1839 = N1837 & N1037;
  assign N1840 = N1838 & N1839;
  assign N1841 = N1840 & N1631;
  assign N1842 = last_r[3] & last_r[2];
  assign N1843 = last_r[1] & N273;
  assign N1844 = N741 & reqs_i[11];
  assign N1845 = N1842 & N1843;
  assign N1846 = N1844 & N1137;
  assign N1847 = N1845 & N1846;
  assign N1848 = N1847 & N349;
  assign N1849 = N1848 & N560;
  assign N1850 = last_r[3] & last_r[2];
  assign N1851 = last_r[1] & N273;
  assign N1852 = N741 & reqs_i[12];
  assign N1853 = N1850 & N1851;
  assign N1854 = N1852 & N1150;
  assign N1855 = N1853 & N1854;
  assign N1856 = N1855 & N447;
  assign N1857 = N1856 & N873;
  assign N1858 = last_r[3] & last_r[2];
  assign N1859 = last_r[1] & N273;
  assign N1860 = N741 & reqs_i[13];
  assign N1861 = N1858 & N1859;
  assign N1862 = N1860 & N1347;
  assign N1863 = N1861 & N1862;
  assign N1864 = N1863 & N544;
  assign N1865 = N1864 & N884;
  assign N1866 = N270 | N271;
  assign N1867 = N272 | last_r[0];
  assign N1868 = reqs_i[15] | N1564;
  assign N1869 = N1866 | N1867;
  assign N1870 = N1868 | N1464;
  assign N1871 = N1869 | N1870;
  assign N1872 = N1871 | N646;
  assign N1873 = N1872 | N1953;
  assign N1875 = last_r[3] & last_r[2];
  assign N1876 = last_r[1] & last_r[0];
  assign N1877 = N1875 & N1876;
  assign N1878 = N1877 & reqs_i[0];
  assign N1879 = last_r[3] & last_r[2];
  assign N1880 = last_r[1] & last_r[0];
  assign N1881 = N1879 & N1880;
  assign N1882 = N1881 & N1476;
  assign N1883 = last_r[3] & last_r[2];
  assign N1884 = last_r[1] & last_r[0];
  assign N1885 = N1883 & N1884;
  assign N1886 = N1885 & N1483;
  assign N1887 = last_r[3] & last_r[2];
  assign N1888 = last_r[1] & last_r[0];
  assign N1889 = N1887 & N1888;
  assign N1890 = N1889 & N1489;
  assign N1891 = last_r[3] & last_r[2];
  assign N1892 = last_r[1] & last_r[0];
  assign N1893 = N1891 & N1892;
  assign N1894 = N1893 & N1495;
  assign N1895 = N1894 & N560;
  assign N1896 = last_r[3] & last_r[2];
  assign N1897 = last_r[1] & last_r[0];
  assign N1898 = N1896 & N1897;
  assign N1899 = N1898 & N400;
  assign N1900 = N1899 & N873;
  assign N1901 = last_r[3] & last_r[2];
  assign N1902 = last_r[1] & last_r[0];
  assign N1903 = N1901 & N1902;
  assign N1904 = N1903 & N497;
  assign N1905 = N1904 & N884;
  assign N1906 = last_r[3] & last_r[2];
  assign N1907 = last_r[1] & last_r[0];
  assign N1908 = N1906 & N1907;
  assign N1909 = N1908 & N595;
  assign N1910 = N1909 & N1598;
  assign N1911 = last_r[3] & last_r[2];
  assign N1912 = last_r[1] & last_r[0];
  assign N1913 = N1911 & N1912;
  assign N1914 = N1913 & N696;
  assign N1915 = N1914 & N1607;
  assign N1916 = last_r[3] & last_r[2];
  assign N1917 = last_r[1] & last_r[0];
  assign N1918 = N1916 & N1917;
  assign N1919 = N1918 & N810;
  assign N1920 = N1919 & N1615;
  assign N1921 = last_r[3] & last_r[2];
  assign N1922 = last_r[1] & last_r[0];
  assign N1923 = N1921 & N1922;
  assign N1924 = N1923 & N916;
  assign N1925 = N1924 & N1623;
  assign N1926 = last_r[3] & last_r[2];
  assign N1927 = last_r[1] & last_r[0];
  assign N1928 = N1926 & N1927;
  assign N1929 = N1928 & N1027;
  assign N1930 = N1929 & N1631;
  assign N1931 = last_r[3] & last_r[2];
  assign N1932 = last_r[1] & last_r[0];
  assign N1933 = N1931 & N1932;
  assign N1934 = N1933 & N1127;
  assign N1935 = N1934 & N349;
  assign N1936 = N1935 & N560;
  assign N1937 = last_r[3] & last_r[2];
  assign N1938 = last_r[1] & last_r[0];
  assign N1939 = N1937 & N1938;
  assign N1940 = N1939 & N1242;
  assign N1941 = N1940 & N447;
  assign N1942 = N1941 & N873;
  assign N1943 = last_r[3] & last_r[2];
  assign N1944 = last_r[1] & last_r[0];
  assign N1945 = N1943 & N1944;
  assign N1946 = N1945 & N1349;
  assign N1947 = N1946 & N544;
  assign N1948 = N1947 & N884;
  assign N1949 = N270 | N271;
  assign N1950 = N272 | N273;
  assign N1951 = reqs_i[1] | reqs_i[0];
  assign N1952 = N1949 | N1950;
  assign N1953 = N457 | N1951;
  assign N1954 = N1952 | N1466;
  assign N1955 = N1954 | N646;
  assign N1956 = N1955 | N1953;
  assign N1958 = N269 | N277 | (N283 | N289) | N296;
  assign N1959 = N303 | N313 | (N319 | N325) | N331;
  assign N1960 = N337 | N344 | (N350 | N356) | N363;
  assign N1961 = N371 | N386 | (N391 | N396) | N401;
  assign N1962 = N406 | N412 | (N418 | N424) | N430;
  assign N1963 = N436 | N442 | (N448 | N454) | N462;
  assign N1964 = N479 | N483 | (N488 | N493) | N498;
  assign N1965 = N503 | N509 | (N515 | N521) | N527;
  assign N1966 = N533 | N539 | (N545 | N552) | N568;
  assign N1967 = N577 | N581 | (N586 | N591) | N596;
  assign N1968 = N601 | N607 | (N613 | N619) | N625;
  assign N1969 = N631 | N637 | (N648 | N661) | N669;
  assign N1970 = N678 | N682 | (N687 | N692) | N697;
  assign N1971 = N702 | N708 | (N714 | N720) | N726;
  assign N1972 = N732 | N740 | (N762 | N772) | N782;
  assign N1973 = N792 | N796 | (N801 | N806) | N811;
  assign N1974 = N816 | N822 | (N828 | N834) | N840;
  assign N1975 = N848 | N862 | (N870 | N879) | N888;
  assign N1976 = N898 | N902 | (N907 | N912) | N917;
  assign N1977 = N923 | N929 | (N935 | N941) | N948;
  assign N1978 = N964 | N972 | (N981 | N990) | N999;
  assign N1979 = N1009 | N1013 | (N1018 | N1023) | N1028;
  assign N1980 = N1034 | N1040 | (N1046 | N1054) | N1066;
  assign N1981 = N1072 | N1078 | (N1085 | N1092) | N1099;
  assign N1982 = N1109 | N1113 | (N1118 | N1123) | N1128;
  assign N1983 = N1134 | N1140 | (N1147 | N1163) | N1171;
  assign N1984 = N1179 | N1187 | (N1196 | N1205) | N1214;
  assign N1985 = N1224 | N1228 | (N1233 | N1238) | N1243;
  assign N1986 = N1249 | N1256 | (N1268 | N1275) | N1282;
  assign N1987 = N1289 | N1296 | (N1304 | N1312) | N1320;
  assign N1988 = N1330 | N1334 | (N1339 | N1344) | N1350;
  assign N1989 = N1356 | N1370 | (N1377 | N1385) | N1393;
  assign N1990 = N1401 | N1409 | (N1418 | N1427) | N1436;
  assign N1991 = N1446 | N1450 | (N1456 | N1461) | N1468;
  assign N1992 = N1479 | N1485 | (N1491 | N1498) | N1504;
  assign N1993 = N1510 | N1516 | (N1523 | N1530) | N1537;
  assign N1994 = N1547 | N1551 | (N1557 | N1563) | N1578;
  assign N1995 = N1585 | N1592 | (N1600 | N1608) | N1616;
  assign N1996 = N1624 | N1632 | (N1640 | N1648) | N1656;
  assign N1997 = N1665 | N1669 | (N1675 | N1685) | N1691;
  assign N1998 = N1697 | N1703 | (N1709 | N1715) | N1721;
  assign N1999 = N1727 | N1733 | (N1740 | N1747) | N1754;
  assign N2000 = N1763 | N1768 | (N1779 | N1785) | N1792;
  assign N2001 = N1799 | N1806 | (N1813 | N1820) | N1827;
  assign N2002 = N1834 | N1841 | (N1849 | N1857) | N1865;
  assign N2003 = N1874 | N1882 | (N1886 | N1890) | N1895;
  assign N2004 = N1900 | N1905 | (N1910 | N1915) | N1920;
  assign N2005 = N1925 | N1930 | (N1936 | N1942) | N1948;
  assign N2006 = N1958 | N1959 | (N1960 | N1961) | N1962;
  assign N2007 = N1963 | N1964 | (N1965 | N1966) | N1967;
  assign N2008 = N1968 | N1969 | (N1970 | N1971) | N1972;
  assign N2009 = N1973 | N1974 | (N1975 | N1976) | N1977;
  assign N2010 = N1978 | N1979 | (N1980 | N1981) | N1982;
  assign N2011 = N1983 | N1984 | (N1985 | N1986) | N1987;
  assign N2012 = N1988 | N1989 | (N1990 | N1991) | N1992;
  assign N2013 = N1993 | N1994 | (N1995 | N1996) | N1997;
  assign N2014 = N1998 | N1999 | (N2000 | N2001) | N2002;
  assign N2015 = N2003 | N2004 | (N2005 | N1957);
  assign N2016 = N2006 | N2007 | (N2008 | N2009) | N2010;
  assign N2017 = N2011 | N2012 | (N2013 | N2014) | N2015;
  assign N2018 = N2016 | N2017;
  assign N2019 = N382 | N470 | (N559 | N654) | N753;
  assign N2020 = N855 | N956 | (N1060 | N1155) | N1262;
  assign N2021 = N1363 | N1473 | (N1571 | N1680) | N1773;
  assign N2022 = N2019 | N2020 | (N2021 | N1878);
  assign N2023 = N269 | N283 | (N289 | N296) | N303;
  assign N2024 = N313 | N319 | (N325 | N331) | N337;
  assign N2025 = N344 | N350 | (N356 | N363) | N371;
  assign N2026 = N382 | N386 | (N391 | N396) | N401;
  assign N2027 = N470 | N483 | (N488 | N493) | N498;
  assign N2028 = N533 | N539 | (N545 | N552) | N559;
  assign N2029 = N631 | N637 | (N648 | N654) | N669;
  assign N2030 = N732 | N740 | (N753 | N772) | N782;
  assign N2031 = N848 | N855 | (N870 | N879) | N888;
  assign N2032 = N956 | N972 | (N981 | N990) | N999;
  assign N2033 = N1034 | N1040 | (N1046 | N1054) | N1060;
  assign N2034 = N1134 | N1140 | (N1147 | N1155) | N1171;
  assign N2035 = N1249 | N1256 | (N1262 | N1275) | N1282;
  assign N2036 = N1356 | N1363 | (N1377 | N1385) | N1393;
  assign N2037 = N1473 | N1485 | (N1491 | N1498) | N1504;
  assign N2038 = N1547 | N1551 | (N1557 | N1563) | N1571;
  assign N2039 = N1665 | N1669 | (N1675 | N1680) | N1691;
  assign N2040 = N1763 | N1768 | (N1773 | N1785) | N1792;
  assign N2041 = N1874 | N1878 | (N1886 | N1890) | N1895;
  assign N2042 = N2023 | N2024 | (N2025 | N2026) | N1962;
  assign N2043 = N1963 | N2027 | (N1965 | N2028) | N1967;
  assign N2044 = N1968 | N2029 | (N1970 | N1971) | N2030;
  assign N2045 = N1973 | N1974 | (N2031 | N1976) | N1977;
  assign N2046 = N2032 | N1979 | (N2033 | N1981) | N1982;
  assign N2047 = N2034 | N1984 | (N1985 | N2035) | N1987;
  assign N2048 = N1988 | N2036 | (N1990 | N1991) | N2037;
  assign N2049 = N1993 | N2038 | (N1995 | N1996) | N2039;
  assign N2050 = N1998 | N1999 | (N2040 | N2001) | N2002;
  assign N2051 = N2041 | N2004 | (N2005 | N1957);
  assign N2052 = N2042 | N2043 | (N2044 | N2045) | N2046;
  assign N2053 = N2047 | N2048 | (N2049 | N2050) | N2051;
  assign N2054 = N2052 | N2053;
  assign N2055 = N277 | N479 | (N568 | N661) | N762;
  assign N2056 = N862 | N964 | (N1066 | N1163) | N1268;
  assign N2057 = N1370 | N1479 | (N1578 | N1685) | N1779;
  assign N2058 = N2055 | N2056 | (N2057 | N1882);
  assign N2059 = N269 | N277 | (N289 | N296) | N303;
  assign N2060 = N382 | N391 | (N396 | N401) | N406;
  assign N2061 = N412 | N418 | (N424 | N430) | N436;
  assign N2062 = N442 | N448 | (N454 | N462) | N470;
  assign N2063 = N568 | N581 | (N586 | N591) | N596;
  assign N2064 = N631 | N637 | (N648 | N654) | N661;
  assign N2065 = N732 | N740 | (N753 | N762) | N782;
  assign N2066 = N848 | N855 | (N862 | N879) | N888;
  assign N2067 = N956 | N964 | (N981 | N990) | N999;
  assign N2068 = N1066 | N1078 | (N1085 | N1092) | N1099;
  assign N2069 = N1134 | N1140 | (N1147 | N1155) | N1163;
  assign N2070 = N1249 | N1256 | (N1262 | N1268) | N1282;
  assign N2071 = N1356 | N1363 | (N1370 | N1385) | N1393;
  assign N2072 = N1473 | N1479 | (N1491 | N1498) | N1504;
  assign N2073 = N1578 | N1592 | (N1600 | N1608) | N1616;
  assign N2074 = N1665 | N1669 | (N1675 | N1680) | N1685;
  assign N2075 = N1763 | N1768 | (N1773 | N1779) | N1792;
  assign N2076 = N1874 | N1878 | (N1882 | N1890) | N1895;
  assign N2077 = N2059 | N2024 | (N2025 | N2060) | N2061;
  assign N2078 = N2062 | N1964 | (N1965 | N2028) | N2063;
  assign N2079 = N1968 | N2064 | (N1970 | N1971) | N2065;
  assign N2080 = N1973 | N1974 | (N2066 | N1976) | N1977;
  assign N2081 = N2067 | N1979 | (N2033 | N2068) | N1982;
  assign N2082 = N2069 | N1984 | (N1985 | N2070) | N1987;
  assign N2083 = N1988 | N2071 | (N1990 | N1991) | N2072;
  assign N2084 = N1993 | N2038 | (N2073 | N1996) | N2074;
  assign N2085 = N1998 | N1999 | (N2075 | N2001) | N2002;
  assign N2086 = N2076 | N2004 | (N2005 | N1957);
  assign N2087 = N2077 | N2078 | (N2079 | N2080) | N2081;
  assign N2088 = N2082 | N2083 | (N2084 | N2085) | N2086;
  assign N2089 = N2087 | N2088;
  assign N2090 = N283 | N386 | (N577 | N669) | N772;
  assign N2091 = N870 | N972 | (N1072 | N1171) | N1275;
  assign N2092 = N1377 | N1485 | (N1585 | N1691) | N1785;
  assign N2093 = N2090 | N2091 | (N2092 | N1886);
  assign N2094 = N269 | N277 | (N283 | N296) | N303;
  assign N2095 = N382 | N386 | (N396 | N401) | N406;
  assign N2096 = N479 | N488 | (N493 | N498) | N503;
  assign N2097 = N509 | N515 | (N521 | N527) | N533;
  assign N2098 = N539 | N545 | (N552 | N559) | N568;
  assign N2099 = N669 | N682 | (N687 | N692) | N697;
  assign N2100 = N732 | N740 | (N753 | N762) | N772;
  assign N2101 = N848 | N855 | (N862 | N870) | N888;
  assign N2102 = N956 | N964 | (N972 | N990) | N999;
  assign N2103 = N1066 | N1072 | (N1085 | N1092) | N1099;
  assign N2104 = N1171 | N1187 | (N1196 | N1205) | N1214;
  assign N2105 = N1249 | N1256 | (N1262 | N1268) | N1275;
  assign N2106 = N1356 | N1363 | (N1370 | N1377) | N1393;
  assign N2107 = N1473 | N1479 | (N1485 | N1498) | N1504;
  assign N2108 = N1578 | N1585 | (N1600 | N1608) | N1616;
  assign N2109 = N1691 | N1703 | (N1709 | N1715) | N1721;
  assign N2110 = N1763 | N1768 | (N1773 | N1779) | N1785;
  assign N2111 = N1874 | N1878 | (N1882 | N1886) | N1895;
  assign N2112 = N2094 | N2024 | (N2025 | N2095) | N2061;
  assign N2113 = N2062 | N2096 | (N2097 | N2098) | N1967;
  assign N2114 = N1968 | N2064 | (N2099 | N1971) | N2100;
  assign N2115 = N1973 | N1974 | (N2101 | N1976) | N1977;
  assign N2116 = N2102 | N1979 | (N2033 | N2103) | N1982;
  assign N2117 = N2069 | N2104 | (N1985 | N2105) | N1987;
  assign N2118 = N1988 | N2106 | (N1990 | N1991) | N2107;
  assign N2119 = N1993 | N2038 | (N2108 | N1996) | N2074;
  assign N2120 = N2109 | N1999 | (N2110 | N2001) | N2002;
  assign N2121 = N2111 | N2004 | (N2005 | N1957);
  assign N2122 = N2112 | N2113 | (N2114 | N2115) | N2116;
  assign N2123 = N2117 | N2118 | (N2119 | N2120) | N2121;
  assign N2124 = N2122 | N2123;
  assign N2125 = N289 | N391 | (N483 | N678) | N782;
  assign N2126 = N879 | N981 | (N1078 | N1179) | N1282;
  assign N2127 = N1385 | N1491 | (N1592 | N1697) | N1792;
  assign N2128 = N2125 | N2126 | (N2127 | N1890);
  assign N2129 = N269 | N277 | (N283 | N289) | N303;
  assign N2130 = N382 | N386 | (N391 | N401) | N406;
  assign N2131 = N479 | N483 | (N493 | N498) | N503;
  assign N2132 = N577 | N586 | (N591 | N596) | N601;
  assign N2133 = N607 | N613 | (N619 | N625) | N631;
  assign N2134 = N637 | N648 | (N654 | N661) | N669;
  assign N2135 = N782 | N796 | (N801 | N806) | N811;
  assign N2136 = N848 | N855 | (N862 | N870) | N879;
  assign N2137 = N956 | N964 | (N972 | N981) | N999;
  assign N2138 = N1066 | N1072 | (N1078 | N1092) | N1099;
  assign N2139 = N1171 | N1179 | (N1196 | N1205) | N1214;
  assign N2140 = N1282 | N1296 | (N1304 | N1312) | N1320;
  assign N2141 = N1356 | N1363 | (N1370 | N1377) | N1385;
  assign N2142 = N1473 | N1479 | (N1485 | N1491) | N1504;
  assign N2143 = N1578 | N1585 | (N1592 | N1608) | N1616;
  assign N2144 = N1691 | N1697 | (N1709 | N1715) | N1721;
  assign N2145 = N1792 | N1806 | (N1813 | N1820) | N1827;
  assign N2146 = N1874 | N1878 | (N1882 | N1886) | N1890;
  assign N2147 = N2129 | N2024 | (N2025 | N2130) | N2061;
  assign N2148 = N2062 | N2131 | (N2097 | N2098) | N2132;
  assign N2149 = N2133 | N2134 | (N1970 | N1971) | N2100;
  assign N2150 = N2135 | N1974 | (N2136 | N1976) | N1977;
  assign N2151 = N2137 | N1979 | (N2033 | N2138) | N1982;
  assign N2152 = N2069 | N2139 | (N1985 | N2105) | N2140;
  assign N2153 = N1988 | N2141 | (N1990 | N1991) | N2142;
  assign N2154 = N1993 | N2038 | (N2143 | N1996) | N2074;
  assign N2155 = N2144 | N1999 | (N2110 | N2145) | N2002;
  assign N2156 = N2146 | N2004 | (N2005 | N1957);
  assign N2157 = N2147 | N2148 | (N2149 | N2150) | N2151;
  assign N2158 = N2152 | N2153 | (N2154 | N2155) | N2156;
  assign N2159 = N2157 | N2158;
  assign N2160 = N296 | N396 | (N488 | N581) | N792;
  assign N2161 = N888 | N990 | (N1085 | N1187) | N1289;
  assign N2162 = N1393 | N1498 | (N1600 | N1703) | N1799;
  assign N2163 = N2160 | N2161 | (N2162 | N1895);
  assign N2164 = N382 | N386 | (N391 | N396) | N406;
  assign N2165 = N479 | N483 | (N488 | N498) | N503;
  assign N2166 = N577 | N581 | (N591 | N596) | N601;
  assign N2167 = N678 | N687 | (N692 | N697) | N702;
  assign N2168 = N708 | N714 | (N720 | N726) | N732;
  assign N2169 = N740 | N753 | (N762 | N772) | N782;
  assign N2170 = N888 | N902 | (N907 | N912) | N917;
  assign N2171 = N956 | N964 | (N972 | N981) | N990;
  assign N2172 = N1066 | N1072 | (N1078 | N1085) | N1099;
  assign N2173 = N1171 | N1179 | (N1187 | N1205) | N1214;
  assign N2174 = N1282 | N1289 | (N1304 | N1312) | N1320;
  assign N2175 = N1393 | N1409 | (N1418 | N1427) | N1436;
  assign N2176 = N1473 | N1479 | (N1485 | N1491) | N1498;
  assign N2177 = N1578 | N1585 | (N1592 | N1600) | N1616;
  assign N2178 = N1691 | N1697 | (N1703 | N1715) | N1721;
  assign N2179 = N1792 | N1799 | (N1813 | N1820) | N1827;
  assign N2180 = N1895 | N1905 | (N1910 | N1915) | N1920;
  assign N2181 = N1958 | N2024 | (N2025 | N2164) | N2061;
  assign N2182 = N2062 | N2165 | (N2097 | N2098) | N2166;
  assign N2183 = N2133 | N2134 | (N2167 | N2168) | N2169;
  assign N2184 = N1973 | N1974 | (N2136 | N2170) | N1977;
  assign N2185 = N2171 | N1979 | (N2033 | N2172) | N1982;
  assign N2186 = N2069 | N2173 | (N1985 | N2105) | N2174;
  assign N2187 = N1988 | N2141 | (N2175 | N1991) | N2176;
  assign N2188 = N1993 | N2038 | (N2177 | N1996) | N2074;
  assign N2189 = N2178 | N1999 | (N2110 | N2179) | N2002;
  assign N2190 = N2146 | N2180 | (N2005 | N1957);
  assign N2191 = N2181 | N2182 | (N2183 | N2184) | N2185;
  assign N2192 = N2186 | N2187 | (N2188 | N2189) | N2190;
  assign N2193 = N2191 | N2192;
  assign N2194 = N303 | N401 | (N493 | N586) | N682;
  assign N2195 = N898 | N999 | (N1092 | N1196) | N1296;
  assign N2196 = N1401 | N1504 | (N1608 | N1709) | N1806;
  assign N2197 = N2194 | N2195 | (N2196 | N1900);
  assign N2198 = N303 | N319 | (N325 | N331) | N337;
  assign N2199 = N479 | N483 | (N488 | N493) | N503;
  assign N2200 = N577 | N581 | (N586 | N596) | N601;
  assign N2201 = N678 | N682 | (N692 | N697) | N702;
  assign N2202 = N792 | N801 | (N806 | N811) | N816;
  assign N2203 = N822 | N828 | (N834 | N840) | N848;
  assign N2204 = N855 | N862 | (N870 | N879) | N888;
  assign N2205 = N999 | N1013 | (N1018 | N1023) | N1028;
  assign N2206 = N1066 | N1072 | (N1078 | N1085) | N1092;
  assign N2207 = N1171 | N1179 | (N1187 | N1196) | N1214;
  assign N2208 = N1282 | N1289 | (N1296 | N1312) | N1320;
  assign N2209 = N1393 | N1401 | (N1418 | N1427) | N1436;
  assign N2210 = N1504 | N1516 | (N1523 | N1530) | N1537;
  assign N2211 = N1578 | N1585 | (N1592 | N1600) | N1608;
  assign N2212 = N1691 | N1697 | (N1703 | N1709) | N1721;
  assign N2213 = N1792 | N1799 | (N1806 | N1820) | N1827;
  assign N2214 = N1895 | N1900 | (N1910 | N1915) | N1920;
  assign N2215 = N1958 | N2198 | (N2025 | N2026) | N2061;
  assign N2216 = N2062 | N2199 | (N2097 | N2098) | N2200;
  assign N2217 = N2133 | N2134 | (N2201 | N2168) | N2169;
  assign N2218 = N2202 | N2203 | (N2204 | N1976) | N1977;
  assign N2219 = N2171 | N2205 | (N2033 | N2206) | N1982;
  assign N2220 = N2069 | N2207 | (N1985 | N2105) | N2208;
  assign N2221 = N1988 | N2141 | (N2209 | N1991) | N2176;
  assign N2222 = N2210 | N2038 | (N2211 | N1996) | N2074;
  assign N2223 = N2212 | N1999 | (N2110 | N2213) | N2002;
  assign N2224 = N2146 | N2214 | (N2005 | N1957);
  assign N2225 = N2215 | N2216 | (N2217 | N2218) | N2219;
  assign N2226 = N2220 | N2221 | (N2222 | N2223) | N2224;
  assign N2227 = N2225 | N2226;
  assign N2228 = N313 | N406 | (N498 | N591) | N687;
  assign N2229 = N796 | N1009 | (N1099 | N1205) | N1304;
  assign N2230 = N1409 | N1510 | (N1616 | N1715) | N1813;
  assign N2231 = N2228 | N2229 | (N2230 | N1905);
  assign N2232 = N303 | N313 | (N325 | N331) | N337;
  assign N2233 = N406 | N418 | (N424 | N430) | N436;
  assign N2234 = N577 | N581 | (N586 | N591) | N601;
  assign N2235 = N678 | N682 | (N687 | N697) | N702;
  assign N2236 = N792 | N796 | (N806 | N811) | N816;
  assign N2237 = N898 | N907 | (N912 | N917) | N923;
  assign N2238 = N929 | N935 | (N941 | N948) | N956;
  assign N2239 = N1099 | N1113 | (N1118 | N1123) | N1128;
  assign N2240 = N1171 | N1179 | (N1187 | N1196) | N1205;
  assign N2241 = N1282 | N1289 | (N1296 | N1304) | N1320;
  assign N2242 = N1393 | N1401 | (N1409 | N1427) | N1436;
  assign N2243 = N1504 | N1510 | (N1523 | N1530) | N1537;
  assign N2244 = N1616 | N1632 | (N1640 | N1648) | N1656;
  assign N2245 = N1691 | N1697 | (N1703 | N1709) | N1715;
  assign N2246 = N1792 | N1799 | (N1806 | N1813) | N1827;
  assign N2247 = N1895 | N1900 | (N1905 | N1915) | N1920;
  assign N2248 = N1958 | N2232 | (N2025 | N2026) | N2233;
  assign N2249 = N2062 | N1964 | (N2097 | N2098) | N2234;
  assign N2250 = N2133 | N2134 | (N2235 | N2168) | N2169;
  assign N2251 = N2236 | N2203 | (N2204 | N2237) | N2238;
  assign N2252 = N1978 | N1979 | (N2033 | N2206) | N2239;
  assign N2253 = N2069 | N2240 | (N1985 | N2105) | N2241;
  assign N2254 = N1988 | N2141 | (N2242 | N1991) | N2176;
  assign N2255 = N2243 | N2038 | (N2211 | N2244) | N2074;
  assign N2256 = N2245 | N1999 | (N2110 | N2246) | N2002;
  assign N2257 = N2146 | N2247 | (N2005 | N1957);
  assign N2258 = N2248 | N2249 | (N2250 | N2251) | N2252;
  assign N2259 = N2253 | N2254 | (N2255 | N2256) | N2257;
  assign N2260 = N2258 | N2259;
  assign N2261 = N319 | N412 | (N503 | N596) | N692;
  assign N2262 = N801 | N902 | (N1109 | N1214) | N1312;
  assign N2263 = N1418 | N1516 | (N1624 | N1721) | N1820;
  assign N2264 = N2261 | N2262 | (N2263 | N1910);
  assign N2265 = N303 | N313 | (N319 | N331) | N337;
  assign N2266 = N406 | N412 | (N424 | N430) | N436;
  assign N2267 = N503 | N515 | (N521 | N527) | N533;
  assign N2268 = N678 | N682 | (N687 | N692) | N702;
  assign N2269 = N792 | N796 | (N801 | N811) | N816;
  assign N2270 = N898 | N902 | (N912 | N917) | N923;
  assign N2271 = N1009 | N1018 | (N1023 | N1028) | N1034;
  assign N2272 = N1040 | N1046 | (N1054 | N1060) | N1066;
  assign N2273 = N1214 | N1228 | (N1233 | N1238) | N1243;
  assign N2274 = N1282 | N1289 | (N1296 | N1304) | N1312;
  assign N2275 = N1393 | N1401 | (N1409 | N1418) | N1436;
  assign N2276 = N1504 | N1510 | (N1516 | N1530) | N1537;
  assign N2277 = N1616 | N1624 | (N1640 | N1648) | N1656;
  assign N2278 = N1721 | N1733 | (N1740 | N1747) | N1754;
  assign N2279 = N1792 | N1799 | (N1806 | N1813) | N1820;
  assign N2280 = N1895 | N1900 | (N1905 | N1910) | N1920;
  assign N2281 = N1958 | N2265 | (N2025 | N2026) | N2266;
  assign N2282 = N2062 | N1964 | (N2267 | N2098) | N1967;
  assign N2283 = N2133 | N2134 | (N2268 | N2168) | N2169;
  assign N2284 = N2269 | N2203 | (N2204 | N2270) | N2238;
  assign N2285 = N1978 | N2271 | (N2272 | N1981) | N1982;
  assign N2286 = N2069 | N2240 | (N2273 | N2105) | N2274;
  assign N2287 = N1988 | N2141 | (N2275 | N1991) | N2176;
  assign N2288 = N2276 | N2038 | (N2211 | N2277) | N2074;
  assign N2289 = N2245 | N2278 | (N2110 | N2279) | N2002;
  assign N2290 = N2146 | N2280 | (N2005 | N1957);
  assign N2291 = N2281 | N2282 | (N2283 | N2284) | N2285;
  assign N2292 = N2286 | N2287 | (N2288 | N2289) | N2290;
  assign N2293 = N2291 | N2292;
  assign N2294 = N325 | N418 | (N509 | N601) | N697;
  assign N2295 = N806 | N907 | (N1013 | N1224) | N1320;
  assign N2296 = N1427 | N1523 | (N1632 | N1727) | N1827;
  assign N2297 = N2294 | N2295 | (N2296 | N1915);
  assign N2298 = N303 | N313 | (N319 | N325) | N337;
  assign N2299 = N406 | N412 | (N418 | N430) | N436;
  assign N2300 = N503 | N509 | (N521 | N527) | N533;
  assign N2301 = N601 | N613 | (N619 | N625) | N631;
  assign N2302 = N792 | N796 | (N801 | N806) | N816;
  assign N2303 = N898 | N902 | (N907 | N917) | N923;
  assign N2304 = N1009 | N1013 | (N1023 | N1028) | N1034;
  assign N2305 = N1109 | N1118 | (N1123 | N1128) | N1134;
  assign N2306 = N1140 | N1147 | (N1155 | N1163) | N1171;
  assign N2307 = N1320 | N1334 | (N1339 | N1344) | N1350;
  assign N2308 = N1393 | N1401 | (N1409 | N1418) | N1427;
  assign N2309 = N1504 | N1510 | (N1516 | N1523) | N1537;
  assign N2310 = N1616 | N1624 | (N1632 | N1648) | N1656;
  assign N2311 = N1721 | N1727 | (N1740 | N1747) | N1754;
  assign N2312 = N1827 | N1841 | (N1849 | N1857) | N1865;
  assign N2313 = N1895 | N1900 | (N1905 | N1910) | N1915;
  assign N2314 = N1958 | N2298 | (N2025 | N2026) | N2299;
  assign N2315 = N2062 | N1964 | (N2300 | N2098) | N1967;
  assign N2316 = N2301 | N2134 | (N1970 | N2168) | N2169;
  assign N2317 = N2302 | N2203 | (N2204 | N2303) | N2238;
  assign N2318 = N1978 | N2304 | (N2272 | N1981) | N2305;
  assign N2319 = N2306 | N1984 | (N1985 | N2105) | N2274;
  assign N2320 = N2307 | N2141 | (N2308 | N1991) | N2176;
  assign N2321 = N2309 | N2038 | (N2211 | N2310) | N2074;
  assign N2322 = N2245 | N2311 | (N2110 | N2279) | N2312;
  assign N2323 = N2146 | N2313 | (N2005 | N1957);
  assign N2324 = N2314 | N2315 | (N2316 | N2317) | N2318;
  assign N2325 = N2319 | N2320 | (N2321 | N2322) | N2323;
  assign N2326 = N2324 | N2325;
  assign N2327 = N331 | N424 | (N515 | N607) | N702;
  assign N2328 = N811 | N912 | (N1018 | N1113) | N1330;
  assign N2329 = N1436 | N1530 | (N1640 | N1733) | N1834;
  assign N2330 = N2327 | N2328 | (N2329 | N1920);
  assign N2331 = N406 | N412 | (N418 | N424) | N436;
  assign N2332 = N503 | N509 | (N515 | N527) | N533;
  assign N2333 = N601 | N607 | (N619 | N625) | N631;
  assign N2334 = N702 | N714 | (N720 | N726) | N732;
  assign N2335 = N898 | N902 | (N907 | N912) | N923;
  assign N2336 = N1009 | N1013 | (N1018 | N1028) | N1034;
  assign N2337 = N1109 | N1113 | (N1123 | N1128) | N1134;
  assign N2338 = N1224 | N1233 | (N1238 | N1243) | N1249;
  assign N2339 = N1256 | N1262 | (N1268 | N1275) | N1282;
  assign N2340 = N1436 | N1450 | (N1456 | N1461) | N1468;
  assign N2341 = N1504 | N1510 | (N1516 | N1523) | N1530;
  assign N2342 = N1616 | N1624 | (N1632 | N1640) | N1656;
  assign N2343 = N1721 | N1727 | (N1733 | N1747) | N1754;
  assign N2344 = N1827 | N1834 | (N1849 | N1857) | N1865;
  assign N2345 = N1920 | N1930 | (N1936 | N1942) | N1948;
  assign N2346 = N1958 | N1959 | (N2025 | N2026) | N2331;
  assign N2347 = N2062 | N1964 | (N2332 | N2098) | N1967;
  assign N2348 = N2333 | N2134 | (N1970 | N2334) | N2169;
  assign N2349 = N1973 | N2203 | (N2204 | N2335) | N2238;
  assign N2350 = N1978 | N2336 | (N2272 | N1981) | N2337;
  assign N2351 = N2306 | N1984 | (N2338 | N2339) | N1987;
  assign N2352 = N1988 | N2141 | (N2308 | N2340) | N2176;
  assign N2353 = N2341 | N2038 | (N2211 | N2342) | N2074;
  assign N2354 = N2245 | N2343 | (N2110 | N2279) | N2344;
  assign N2355 = N2146 | N2313 | (N2345 | N1957);
  assign N2356 = N2346 | N2347 | (N2348 | N2349) | N2350;
  assign N2357 = N2351 | N2352 | (N2353 | N2354) | N2355;
  assign N2358 = N2356 | N2357;
  assign N2359 = N337 | N430 | (N521 | N613) | N708;
  assign N2360 = N816 | N917 | (N1023 | N1118) | N1228;
  assign N2361 = N1446 | N1537 | (N1648 | N1740) | N1841;
  assign N2362 = N2359 | N2360 | (N2361 | N1925);
  assign N2363 = N337 | N350 | (N356 | N363) | N371;
  assign N2364 = N503 | N509 | (N515 | N521) | N533;
  assign N2365 = N601 | N607 | (N613 | N625) | N631;
  assign N2366 = N702 | N708 | (N720 | N726) | N732;
  assign N2367 = N816 | N828 | (N834 | N840) | N848;
  assign N2368 = N1009 | N1013 | (N1018 | N1023) | N1034;
  assign N2369 = N1109 | N1113 | (N1118 | N1128) | N1134;
  assign N2370 = N1224 | N1228 | (N1238 | N1243) | N1249;
  assign N2371 = N1330 | N1339 | (N1344 | N1350) | N1356;
  assign N2372 = N1363 | N1370 | (N1377 | N1385) | N1393;
  assign N2373 = N1537 | N1551 | (N1557 | N1563) | N1571;
  assign N2374 = N1616 | N1624 | (N1632 | N1640) | N1648;
  assign N2375 = N1721 | N1727 | (N1733 | N1740) | N1754;
  assign N2376 = N1827 | N1834 | (N1841 | N1857) | N1865;
  assign N2377 = N1920 | N1925 | (N1936 | N1942) | N1948;
  assign N2378 = N1958 | N1959 | (N2363 | N2026) | N1962;
  assign N2379 = N2062 | N1964 | (N2364 | N2098) | N1967;
  assign N2380 = N2365 | N2134 | (N1970 | N2366) | N2169;
  assign N2381 = N1973 | N2367 | (N2204 | N1976) | N2238;
  assign N2382 = N1978 | N2368 | (N2272 | N1981) | N2369;
  assign N2383 = N2306 | N1984 | (N2370 | N2339) | N1987;
  assign N2384 = N2371 | N2372 | (N1990 | N1991) | N2176;
  assign N2385 = N2341 | N2373 | (N2211 | N2374) | N2074;
  assign N2386 = N2245 | N2375 | (N2110 | N2279) | N2376;
  assign N2387 = N2146 | N2313 | (N2377 | N1957);
  assign N2388 = N2378 | N2379 | (N2380 | N2381) | N2382;
  assign N2389 = N2383 | N2384 | (N2385 | N2386) | N2387;
  assign N2390 = N2388 | N2389;
  assign N2391 = N344 | N436 | (N527 | N619) | N714;
  assign N2392 = N822 | N923 | (N1028 | N1123) | N1233;
  assign N2393 = N1334 | N1547 | (N1656 | N1747) | N1849;
  assign N2394 = N2391 | N2392 | (N2393 | N1930);
  assign N2395 = N337 | N344 | (N356 | N363) | N371;
  assign N2396 = N436 | N448 | (N454 | N462) | N470;
  assign N2397 = N601 | N607 | (N613 | N619) | N631;
  assign N2398 = N702 | N708 | (N714 | N726) | N732;
  assign N2399 = N816 | N822 | (N834 | N840) | N848;
  assign N2400 = N923 | N935 | (N941 | N948) | N956;
  assign N2401 = N1109 | N1113 | (N1118 | N1123) | N1134;
  assign N2402 = N1224 | N1228 | (N1233 | N1243) | N1249;
  assign N2403 = N1330 | N1334 | (N1344 | N1350) | N1356;
  assign N2404 = N1446 | N1456 | (N1461 | N1468) | N1473;
  assign N2405 = N1656 | N1669 | (N1675 | N1680) | N1685;
  assign N2406 = N1721 | N1727 | (N1733 | N1740) | N1747;
  assign N2407 = N1827 | N1834 | (N1841 | N1849) | N1865;
  assign N2408 = N1920 | N1925 | (N1930 | N1942) | N1948;
  assign N2409 = N1958 | N1959 | (N2395 | N2026) | N1962;
  assign N2410 = N2396 | N1964 | (N1965 | N2098) | N1967;
  assign N2411 = N2397 | N2134 | (N1970 | N2398) | N2169;
  assign N2412 = N1973 | N2399 | (N2204 | N1976) | N2400;
  assign N2413 = N1978 | N1979 | (N2272 | N1981) | N2401;
  assign N2414 = N2306 | N1984 | (N2402 | N2339) | N1987;
  assign N2415 = N2403 | N2372 | (N1990 | N2404) | N1992;
  assign N2416 = N1993 | N2038 | (N2211 | N2374) | N2405;
  assign N2417 = N2245 | N2406 | (N2110 | N2279) | N2407;
  assign N2418 = N2146 | N2313 | (N2408 | N1957);
  assign N2419 = N2409 | N2410 | (N2411 | N2412) | N2413;
  assign N2420 = N2414 | N2415 | (N2416 | N2417) | N2418;
  assign N2421 = N2419 | N2420;
  assign N2422 = N350 | N442 | (N533 | N625) | N720;
  assign N2423 = N828 | N929 | (N1034 | N1128) | N1238;
  assign N2424 = N1339 | N1450 | (N1665 | N1754) | N1857;
  assign N2425 = N2422 | N2423 | (N2424 | N1936);
  assign N2426 = N337 | N344 | (N350 | N363) | N371;
  assign N2427 = N436 | N442 | (N454 | N462) | N470;
  assign N2428 = N533 | N545 | (N552 | N559) | N568;
  assign N2429 = N702 | N708 | (N714 | N720) | N732;
  assign N2430 = N816 | N822 | (N828 | N840) | N848;
  assign N2431 = N923 | N929 | (N941 | N948) | N956;
  assign N2432 = N1034 | N1046 | (N1054 | N1060) | N1066;
  assign N2433 = N1224 | N1228 | (N1233 | N1238) | N1249;
  assign N2434 = N1330 | N1334 | (N1339 | N1350) | N1356;
  assign N2435 = N1446 | N1450 | (N1461 | N1468) | N1473;
  assign N2436 = N1547 | N1557 | (N1563 | N1571) | N1578;
  assign N2437 = N1754 | N1768 | (N1773 | N1779) | N1785;
  assign N2438 = N1827 | N1834 | (N1841 | N1849) | N1857;
  assign N2439 = N1920 | N1925 | (N1930 | N1936) | N1948;
  assign N2440 = N1958 | N1959 | (N2426 | N2026) | N1962;
  assign N2441 = N2427 | N1964 | (N1965 | N2428) | N1967;
  assign N2442 = N1968 | N2134 | (N1970 | N2429) | N2169;
  assign N2443 = N1973 | N2430 | (N2204 | N1976) | N2431;
  assign N2444 = N1978 | N1979 | (N2432 | N1981) | N1982;
  assign N2445 = N2306 | N1984 | (N2433 | N2339) | N1987;
  assign N2446 = N2434 | N2372 | (N1990 | N2435) | N1992;
  assign N2447 = N1993 | N2436 | (N1995 | N1996) | N2074;
  assign N2448 = N2245 | N2406 | (N2437 | N2279) | N2438;
  assign N2449 = N2146 | N2313 | (N2439 | N1957);
  assign N2450 = N2440 | N2441 | (N2442 | N2443) | N2444;
  assign N2451 = N2445 | N2446 | (N2447 | N2448) | N2449;
  assign N2452 = N2450 | N2451;
  assign N2453 = N356 | N448 | (N539 | N631) | N726;
  assign N2454 = N834 | N935 | (N1040 | N1134) | N1243;
  assign N2455 = N1344 | N1456 | (N1551 | N1763) | N1865;
  assign N2456 = N2453 | N2454 | (N2455 | N1942);
  assign N2457 = N337 | N344 | (N350 | N356) | N371;
  assign N2458 = N436 | N442 | (N448 | N462) | N470;
  assign N2459 = N533 | N539 | (N552 | N559) | N568;
  assign N2460 = N631 | N648 | (N654 | N661) | N669;
  assign N2461 = N816 | N822 | (N828 | N834) | N848;
  assign N2462 = N923 | N929 | (N935 | N948) | N956;
  assign N2463 = N1034 | N1040 | (N1054 | N1060) | N1066;
  assign N2464 = N1134 | N1147 | (N1155 | N1163) | N1171;
  assign N2465 = N1330 | N1334 | (N1339 | N1344) | N1356;
  assign N2466 = N1446 | N1450 | (N1456 | N1468) | N1473;
  assign N2467 = N1547 | N1551 | (N1563 | N1571) | N1578;
  assign N2468 = N1665 | N1675 | (N1680 | N1685) | N1691;
  assign N2469 = N1865 | N1878 | (N1882 | N1886) | N1890;
  assign N2470 = N1920 | N1925 | (N1930 | N1936) | N1942;
  assign N2471 = N1958 | N1959 | (N2457 | N2026) | N1962;
  assign N2472 = N2458 | N1964 | (N1965 | N2459) | N1967;
  assign N2473 = N1968 | N2460 | (N1970 | N1971) | N2169;
  assign N2474 = N1973 | N2461 | (N2204 | N1976) | N2462;
  assign N2475 = N1978 | N1979 | (N2463 | N1981) | N1982;
  assign N2476 = N2464 | N1984 | (N1985 | N2339) | N1987;
  assign N2477 = N2465 | N2372 | (N1990 | N2466) | N1992;
  assign N2478 = N1993 | N2467 | (N1995 | N1996) | N2468;
  assign N2479 = N1998 | N1999 | (N2110 | N2279) | N2438;
  assign N2480 = N2469 | N2313 | (N2470 | N1957);
  assign N2481 = N2471 | N2472 | (N2473 | N2474) | N2475;
  assign N2482 = N2476 | N2477 | (N2478 | N2479) | N2480;
  assign N2483 = N2481 | N2482;
  assign N2484 = N363 | N454 | (N545 | N637) | N732;
  assign N2485 = N840 | N941 | (N1046 | N1140) | N1249;
  assign N2486 = N1350 | N1461 | (N1557 | N1669) | N1874;
  assign N2487 = N2484 | N2485 | (N2486 | N1948);
  assign N2488 = N436 | N442 | (N448 | N454) | N470;
  assign N2489 = N533 | N539 | (N545 | N559) | N568;
  assign N2490 = N631 | N637 | (N654 | N661) | N669;
  assign N2491 = N732 | N753 | (N762 | N772) | N782;
  assign N2492 = N923 | N929 | (N935 | N941) | N956;
  assign N2493 = N1034 | N1040 | (N1046 | N1060) | N1066;
  assign N2494 = N1134 | N1140 | (N1155 | N1163) | N1171;
  assign N2495 = N1249 | N1262 | (N1268 | N1275) | N1282;
  assign N2496 = N1446 | N1450 | (N1456 | N1461) | N1473;
  assign N2497 = N1547 | N1551 | (N1557 | N1571) | N1578;
  assign N2498 = N1665 | N1669 | (N1680 | N1685) | N1691;
  assign N2499 = N1763 | N1773 | (N1779 | N1785) | N1792;
  assign N2500 = N1958 | N1959 | (N1960 | N2026) | N1962;
  assign N2501 = N2488 | N1964 | (N1965 | N2489) | N1967;
  assign N2502 = N1968 | N2490 | (N1970 | N1971) | N2491;
  assign N2503 = N1973 | N1974 | (N2204 | N1976) | N2492;
  assign N2504 = N1978 | N1979 | (N2493 | N1981) | N1982;
  assign N2505 = N2494 | N1984 | (N1985 | N2495) | N1987;
  assign N2506 = N1988 | N2372 | (N1990 | N2496) | N1992;
  assign N2507 = N1993 | N2497 | (N1995 | N1996) | N2498;
  assign N2508 = N1998 | N1999 | (N2499 | N2001) | N2002;
  assign N2509 = N2146 | N2313 | (N2470 | N1948);
  assign N2510 = N2500 | N2501 | (N2502 | N2503) | N2504;
  assign N2511 = N2505 | N2506 | (N2507 | N2508) | N2509;
  assign N2512 = N2510 | N2511;
  assign N2513 = N371 | N462 | (N552 | N648) | N740;
  assign N2514 = N848 | N948 | (N1054 | N1147) | N1256;
  assign N2515 = N1356 | N1468 | (N1563 | N1675) | N1768;
  assign N2516 = N2513 | N2514 | (N2515 | N1957);
  assign sel_one_hot_o[0] = (N0)? 1'b0 : 
                            (N1)? 1'b1 : 1'b0;
  assign N0 = N2018;
  assign N1 = N2022;
  assign sel_one_hot_o[1] = (N2)? 1'b0 : 
                            (N3)? 1'b1 : 1'b0;
  assign N2 = N2054;
  assign N3 = N2058;
  assign sel_one_hot_o[2] = (N4)? 1'b0 : 
                            (N5)? 1'b1 : 1'b0;
  assign N4 = N2089;
  assign N5 = N2093;
  assign sel_one_hot_o[3] = (N6)? 1'b0 : 
                            (N7)? 1'b1 : 1'b0;
  assign N6 = N2124;
  assign N7 = N2128;
  assign sel_one_hot_o[4] = (N8)? 1'b0 : 
                            (N9)? 1'b1 : 1'b0;
  assign N8 = N2159;
  assign N9 = N2163;
  assign sel_one_hot_o[5] = (N10)? 1'b0 : 
                            (N11)? 1'b1 : 1'b0;
  assign N10 = N2193;
  assign N11 = N2197;
  assign sel_one_hot_o[6] = (N12)? 1'b0 : 
                            (N13)? 1'b1 : 1'b0;
  assign N12 = N2227;
  assign N13 = N2231;
  assign sel_one_hot_o[7] = (N14)? 1'b0 : 
                            (N15)? 1'b1 : 1'b0;
  assign N14 = N2260;
  assign N15 = N2264;
  assign sel_one_hot_o[8] = (N16)? 1'b0 : 
                            (N17)? 1'b1 : 1'b0;
  assign N16 = N2293;
  assign N17 = N2297;
  assign sel_one_hot_o[9] = (N18)? 1'b0 : 
                            (N19)? 1'b1 : 1'b0;
  assign N18 = N2326;
  assign N19 = N2330;
  assign sel_one_hot_o[10] = (N20)? 1'b0 : 
                             (N21)? 1'b1 : 1'b0;
  assign N20 = N2358;
  assign N21 = N2362;
  assign sel_one_hot_o[11] = (N22)? 1'b0 : 
                             (N23)? 1'b1 : 1'b0;
  assign N22 = N2390;
  assign N23 = N2394;
  assign sel_one_hot_o[12] = (N24)? 1'b0 : 
                             (N25)? 1'b1 : 1'b0;
  assign N24 = N2421;
  assign N25 = N2425;
  assign sel_one_hot_o[13] = (N26)? 1'b0 : 
                             (N27)? 1'b1 : 1'b0;
  assign N26 = N2452;
  assign N27 = N2456;
  assign sel_one_hot_o[14] = (N28)? 1'b0 : 
                             (N29)? 1'b1 : 1'b0;
  assign N28 = N2483;
  assign N29 = N2487;
  assign sel_one_hot_o[15] = (N30)? 1'b0 : 
                             (N31)? 1'b1 : 1'b0;
  assign N30 = N2512;
  assign N31 = N2516;
  assign tag_o[3] = (N32)? 1'b0 : 
                    (N33)? 1'b0 : 
                    (N34)? 1'b0 : 
                    (N35)? 1'b0 : 
                    (N36)? 1'b0 : 
                    (N37)? 1'b0 : 
                    (N38)? 1'b0 : 
                    (N39)? 1'b0 : 
                    (N40)? 1'b1 : 
                    (N41)? 1'b1 : 
                    (N42)? 1'b1 : 
                    (N43)? 1'b1 : 
                    (N44)? 1'b1 : 
                    (N45)? 1'b1 : 
                    (N46)? 1'b1 : 
                    (N371)? 1'b1 : 
                    (N382)? 1'b0 : 
                    (N47)? 1'b0 : 
                    (N48)? 1'b0 : 
                    (N49)? 1'b0 : 
                    (N50)? 1'b0 : 
                    (N51)? 1'b0 : 
                    (N52)? 1'b0 : 
                    (N53)? 1'b1 : 
                    (N54)? 1'b1 : 
                    (N55)? 1'b1 : 
                    (N56)? 1'b1 : 
                    (N57)? 1'b1 : 
                    (N58)? 1'b1 : 
                    (N59)? 1'b1 : 
                    (N462)? 1'b1 : 
                    (N60)? 1'b0 : 
                    (N479)? 1'b0 : 
                    (N61)? 1'b0 : 
                    (N62)? 1'b0 : 
                    (N63)? 1'b0 : 
                    (N64)? 1'b0 : 
                    (N65)? 1'b0 : 
                    (N66)? 1'b1 : 
                    (N67)? 1'b1 : 
                    (N68)? 1'b1 : 
                    (N69)? 1'b1 : 
                    (N70)? 1'b1 : 
                    (N71)? 1'b1 : 
                    (N72)? 1'b1 : 
                    (N552)? 1'b1 : 
                    (N73)? 1'b0 : 
                    (N74)? 1'b0 : 
                    (N577)? 1'b0 : 
                    (N75)? 1'b0 : 
                    (N76)? 1'b0 : 
                    (N77)? 1'b0 : 
                    (N78)? 1'b0 : 
                    (N79)? 1'b1 : 
                    (N80)? 1'b1 : 
                    (N81)? 1'b1 : 
                    (N82)? 1'b1 : 
                    (N83)? 1'b1 : 
                    (N84)? 1'b1 : 
                    (N85)? 1'b1 : 
                    (N648)? 1'b1 : 
                    (N86)? 1'b0 : 
                    (N87)? 1'b0 : 
                    (N88)? 1'b0 : 
                    (N678)? 1'b0 : 
                    (N89)? 1'b0 : 
                    (N90)? 1'b0 : 
                    (N91)? 1'b0 : 
                    (N92)? 1'b1 : 
                    (N93)? 1'b1 : 
                    (N94)? 1'b1 : 
                    (N95)? 1'b1 : 
                    (N96)? 1'b1 : 
                    (N97)? 1'b1 : 
                    (N98)? 1'b1 : 
                    (N740)? 1'b1 : 
                    (N99)? 1'b0 : 
                    (N100)? 1'b0 : 
                    (N101)? 1'b0 : 
                    (N102)? 1'b0 : 
                    (N792)? 1'b0 : 
                    (N103)? 1'b0 : 
                    (N104)? 1'b0 : 
                    (N105)? 1'b1 : 
                    (N106)? 1'b1 : 
                    (N107)? 1'b1 : 
                    (N108)? 1'b1 : 
                    (N109)? 1'b1 : 
                    (N110)? 1'b1 : 
                    (N111)? 1'b1 : 
                    (N848)? 1'b1 : 
                    (N112)? 1'b0 : 
                    (N113)? 1'b0 : 
                    (N114)? 1'b0 : 
                    (N115)? 1'b0 : 
                    (N116)? 1'b0 : 
                    (N898)? 1'b0 : 
                    (N117)? 1'b0 : 
                    (N118)? 1'b1 : 
                    (N119)? 1'b1 : 
                    (N120)? 1'b1 : 
                    (N121)? 1'b1 : 
                    (N122)? 1'b1 : 
                    (N123)? 1'b1 : 
                    (N124)? 1'b1 : 
                    (N948)? 1'b1 : 
                    (N125)? 1'b0 : 
                    (N126)? 1'b0 : 
                    (N127)? 1'b0 : 
                    (N128)? 1'b0 : 
                    (N129)? 1'b0 : 
                    (N130)? 1'b0 : 
                    (N1009)? 1'b0 : 
                    (N131)? 1'b1 : 
                    (N132)? 1'b1 : 
                    (N133)? 1'b1 : 
                    (N134)? 1'b1 : 
                    (N135)? 1'b1 : 
                    (N136)? 1'b1 : 
                    (N137)? 1'b1 : 
                    (N1054)? 1'b1 : 
                    (N138)? 1'b0 : 
                    (N139)? 1'b0 : 
                    (N140)? 1'b0 : 
                    (N141)? 1'b0 : 
                    (N142)? 1'b0 : 
                    (N143)? 1'b0 : 
                    (N144)? 1'b0 : 
                    (N1109)? 1'b0 : 
                    (N145)? 1'b1 : 
                    (N146)? 1'b1 : 
                    (N147)? 1'b1 : 
                    (N148)? 1'b1 : 
                    (N149)? 1'b1 : 
                    (N150)? 1'b1 : 
                    (N1147)? 1'b1 : 
                    (N151)? 1'b0 : 
                    (N152)? 1'b0 : 
                    (N153)? 1'b0 : 
                    (N154)? 1'b0 : 
                    (N155)? 1'b0 : 
                    (N156)? 1'b0 : 
                    (N157)? 1'b0 : 
                    (N158)? 1'b0 : 
                    (N1224)? 1'b1 : 
                    (N159)? 1'b1 : 
                    (N160)? 1'b1 : 
                    (N161)? 1'b1 : 
                    (N162)? 1'b1 : 
                    (N163)? 1'b1 : 
                    (N1256)? 1'b1 : 
                    (N164)? 1'b0 : 
                    (N165)? 1'b0 : 
                    (N166)? 1'b0 : 
                    (N167)? 1'b0 : 
                    (N168)? 1'b0 : 
                    (N169)? 1'b0 : 
                    (N170)? 1'b0 : 
                    (N171)? 1'b0 : 
                    (N172)? 1'b1 : 
                    (N1330)? 1'b1 : 
                    (N173)? 1'b1 : 
                    (N174)? 1'b1 : 
                    (N175)? 1'b1 : 
                    (N176)? 1'b1 : 
                    (N1356)? 1'b1 : 
                    (N177)? 1'b0 : 
                    (N178)? 1'b0 : 
                    (N179)? 1'b0 : 
                    (N180)? 1'b0 : 
                    (N181)? 1'b0 : 
                    (N182)? 1'b0 : 
                    (N183)? 1'b0 : 
                    (N184)? 1'b0 : 
                    (N185)? 1'b1 : 
                    (N186)? 1'b1 : 
                    (N1446)? 1'b1 : 
                    (N187)? 1'b1 : 
                    (N188)? 1'b1 : 
                    (N189)? 1'b1 : 
                    (N1468)? 1'b1 : 
                    (N190)? 1'b0 : 
                    (N191)? 1'b0 : 
                    (N192)? 1'b0 : 
                    (N193)? 1'b0 : 
                    (N194)? 1'b0 : 
                    (N195)? 1'b0 : 
                    (N196)? 1'b0 : 
                    (N197)? 1'b0 : 
                    (N198)? 1'b1 : 
                    (N199)? 1'b1 : 
                    (N200)? 1'b1 : 
                    (N1547)? 1'b1 : 
                    (N201)? 1'b1 : 
                    (N202)? 1'b1 : 
                    (N1563)? 1'b1 : 
                    (N203)? 1'b0 : 
                    (N204)? 1'b0 : 
                    (N205)? 1'b0 : 
                    (N206)? 1'b0 : 
                    (N207)? 1'b0 : 
                    (N208)? 1'b0 : 
                    (N209)? 1'b0 : 
                    (N210)? 1'b0 : 
                    (N211)? 1'b1 : 
                    (N212)? 1'b1 : 
                    (N213)? 1'b1 : 
                    (N214)? 1'b1 : 
                    (N1665)? 1'b1 : 
                    (N215)? 1'b1 : 
                    (N1675)? 1'b1 : 
                    (N216)? 1'b0 : 
                    (N217)? 1'b0 : 
                    (N218)? 1'b0 : 
                    (N219)? 1'b0 : 
                    (N220)? 1'b0 : 
                    (N221)? 1'b0 : 
                    (N222)? 1'b0 : 
                    (N223)? 1'b0 : 
                    (N224)? 1'b1 : 
                    (N225)? 1'b1 : 
                    (N226)? 1'b1 : 
                    (N227)? 1'b1 : 
                    (N228)? 1'b1 : 
                    (N1763)? 1'b1 : 
                    (N1768)? 1'b1 : 
                    (N229)? 1'b0 : 
                    (N230)? 1'b0 : 
                    (N231)? 1'b0 : 
                    (N232)? 1'b0 : 
                    (N233)? 1'b0 : 
                    (N234)? 1'b0 : 
                    (N235)? 1'b0 : 
                    (N236)? 1'b0 : 
                    (N237)? 1'b1 : 
                    (N238)? 1'b1 : 
                    (N239)? 1'b1 : 
                    (N240)? 1'b1 : 
                    (N241)? 1'b1 : 
                    (N242)? 1'b1 : 
                    (N1874)? 1'b1 : 
                    (N243)? 1'b0 : 
                    (N244)? 1'b0 : 
                    (N245)? 1'b0 : 
                    (N246)? 1'b0 : 
                    (N247)? 1'b0 : 
                    (N248)? 1'b0 : 
                    (N249)? 1'b0 : 
                    (N250)? 1'b0 : 
                    (N251)? 1'b1 : 
                    (N252)? 1'b1 : 
                    (N253)? 1'b1 : 
                    (N254)? 1'b1 : 
                    (N255)? 1'b1 : 
                    (N256)? 1'b1 : 
                    (N257)? 1'b1 : 
                    (N1957)? 1'b1 : 1'b0;
  assign N32 = N269;
  assign N33 = N277;
  assign N34 = N283;
  assign N35 = N289;
  assign N36 = N296;
  assign N37 = N303;
  assign N38 = N313;
  assign N39 = N319;
  assign N40 = N325;
  assign N41 = N331;
  assign N42 = N337;
  assign N43 = N344;
  assign N44 = N350;
  assign N45 = N356;
  assign N46 = N363;
  assign N47 = N386;
  assign N48 = N391;
  assign N49 = N396;
  assign N50 = N401;
  assign N51 = N406;
  assign N52 = N412;
  assign N53 = N418;
  assign N54 = N424;
  assign N55 = N430;
  assign N56 = N436;
  assign N57 = N442;
  assign N58 = N448;
  assign N59 = N454;
  assign N60 = N470;
  assign N61 = N483;
  assign N62 = N488;
  assign N63 = N493;
  assign N64 = N498;
  assign N65 = N503;
  assign N66 = N509;
  assign N67 = N515;
  assign N68 = N521;
  assign N69 = N527;
  assign N70 = N533;
  assign N71 = N539;
  assign N72 = N545;
  assign N73 = N559;
  assign N74 = N568;
  assign N75 = N581;
  assign N76 = N586;
  assign N77 = N591;
  assign N78 = N596;
  assign N79 = N601;
  assign N80 = N607;
  assign N81 = N613;
  assign N82 = N619;
  assign N83 = N625;
  assign N84 = N631;
  assign N85 = N637;
  assign N86 = N654;
  assign N87 = N661;
  assign N88 = N669;
  assign N89 = N682;
  assign N90 = N687;
  assign N91 = N692;
  assign N92 = N697;
  assign N93 = N702;
  assign N94 = N708;
  assign N95 = N714;
  assign N96 = N720;
  assign N97 = N726;
  assign N98 = N732;
  assign N99 = N753;
  assign N100 = N762;
  assign N101 = N772;
  assign N102 = N782;
  assign N103 = N796;
  assign N104 = N801;
  assign N105 = N806;
  assign N106 = N811;
  assign N107 = N816;
  assign N108 = N822;
  assign N109 = N828;
  assign N110 = N834;
  assign N111 = N840;
  assign N112 = N855;
  assign N113 = N862;
  assign N114 = N870;
  assign N115 = N879;
  assign N116 = N888;
  assign N117 = N902;
  assign N118 = N907;
  assign N119 = N912;
  assign N120 = N917;
  assign N121 = N923;
  assign N122 = N929;
  assign N123 = N935;
  assign N124 = N941;
  assign N125 = N956;
  assign N126 = N964;
  assign N127 = N972;
  assign N128 = N981;
  assign N129 = N990;
  assign N130 = N999;
  assign N131 = N1013;
  assign N132 = N1018;
  assign N133 = N1023;
  assign N134 = N1028;
  assign N135 = N1034;
  assign N136 = N1040;
  assign N137 = N1046;
  assign N138 = N1060;
  assign N139 = N1066;
  assign N140 = N1072;
  assign N141 = N1078;
  assign N142 = N1085;
  assign N143 = N1092;
  assign N144 = N1099;
  assign N145 = N1113;
  assign N146 = N1118;
  assign N147 = N1123;
  assign N148 = N1128;
  assign N149 = N1134;
  assign N150 = N1140;
  assign N151 = N1155;
  assign N152 = N1163;
  assign N153 = N1171;
  assign N154 = N1179;
  assign N155 = N1187;
  assign N156 = N1196;
  assign N157 = N1205;
  assign N158 = N1214;
  assign N159 = N1228;
  assign N160 = N1233;
  assign N161 = N1238;
  assign N162 = N1243;
  assign N163 = N1249;
  assign N164 = N1262;
  assign N165 = N1268;
  assign N166 = N1275;
  assign N167 = N1282;
  assign N168 = N1289;
  assign N169 = N1296;
  assign N170 = N1304;
  assign N171 = N1312;
  assign N172 = N1320;
  assign N173 = N1334;
  assign N174 = N1339;
  assign N175 = N1344;
  assign N176 = N1350;
  assign N177 = N1363;
  assign N178 = N1370;
  assign N179 = N1377;
  assign N180 = N1385;
  assign N181 = N1393;
  assign N182 = N1401;
  assign N183 = N1409;
  assign N184 = N1418;
  assign N185 = N1427;
  assign N186 = N1436;
  assign N187 = N1450;
  assign N188 = N1456;
  assign N189 = N1461;
  assign N190 = N1473;
  assign N191 = N1479;
  assign N192 = N1485;
  assign N193 = N1491;
  assign N194 = N1498;
  assign N195 = N1504;
  assign N196 = N1510;
  assign N197 = N1516;
  assign N198 = N1523;
  assign N199 = N1530;
  assign N200 = N1537;
  assign N201 = N1551;
  assign N202 = N1557;
  assign N203 = N1571;
  assign N204 = N1578;
  assign N205 = N1585;
  assign N206 = N1592;
  assign N207 = N1600;
  assign N208 = N1608;
  assign N209 = N1616;
  assign N210 = N1624;
  assign N211 = N1632;
  assign N212 = N1640;
  assign N213 = N1648;
  assign N214 = N1656;
  assign N215 = N1669;
  assign N216 = N1680;
  assign N217 = N1685;
  assign N218 = N1691;
  assign N219 = N1697;
  assign N220 = N1703;
  assign N221 = N1709;
  assign N222 = N1715;
  assign N223 = N1721;
  assign N224 = N1727;
  assign N225 = N1733;
  assign N226 = N1740;
  assign N227 = N1747;
  assign N228 = N1754;
  assign N229 = N1773;
  assign N230 = N1779;
  assign N231 = N1785;
  assign N232 = N1792;
  assign N233 = N1799;
  assign N234 = N1806;
  assign N235 = N1813;
  assign N236 = N1820;
  assign N237 = N1827;
  assign N238 = N1834;
  assign N239 = N1841;
  assign N240 = N1849;
  assign N241 = N1857;
  assign N242 = N1865;
  assign N243 = N1878;
  assign N244 = N1882;
  assign N245 = N1886;
  assign N246 = N1890;
  assign N247 = N1895;
  assign N248 = N1900;
  assign N249 = N1905;
  assign N250 = N1910;
  assign N251 = N1915;
  assign N252 = N1920;
  assign N253 = N1925;
  assign N254 = N1930;
  assign N255 = N1936;
  assign N256 = N1942;
  assign N257 = N1948;
  assign tag_o[2] = (N32)? 1'b0 : 
                    (N33)? 1'b0 : 
                    (N34)? 1'b0 : 
                    (N35)? 1'b0 : 
                    (N36)? 1'b1 : 
                    (N37)? 1'b1 : 
                    (N38)? 1'b1 : 
                    (N39)? 1'b1 : 
                    (N40)? 1'b0 : 
                    (N41)? 1'b0 : 
                    (N42)? 1'b0 : 
                    (N43)? 1'b0 : 
                    (N44)? 1'b1 : 
                    (N45)? 1'b1 : 
                    (N46)? 1'b1 : 
                    (N371)? 1'b1 : 
                    (N382)? 1'b0 : 
                    (N47)? 1'b0 : 
                    (N48)? 1'b0 : 
                    (N49)? 1'b1 : 
                    (N50)? 1'b1 : 
                    (N51)? 1'b1 : 
                    (N52)? 1'b1 : 
                    (N53)? 1'b0 : 
                    (N54)? 1'b0 : 
                    (N55)? 1'b0 : 
                    (N56)? 1'b0 : 
                    (N57)? 1'b1 : 
                    (N58)? 1'b1 : 
                    (N59)? 1'b1 : 
                    (N462)? 1'b1 : 
                    (N60)? 1'b0 : 
                    (N479)? 1'b0 : 
                    (N61)? 1'b0 : 
                    (N62)? 1'b1 : 
                    (N63)? 1'b1 : 
                    (N64)? 1'b1 : 
                    (N65)? 1'b1 : 
                    (N66)? 1'b0 : 
                    (N67)? 1'b0 : 
                    (N68)? 1'b0 : 
                    (N69)? 1'b0 : 
                    (N70)? 1'b1 : 
                    (N71)? 1'b1 : 
                    (N72)? 1'b1 : 
                    (N552)? 1'b1 : 
                    (N73)? 1'b0 : 
                    (N74)? 1'b0 : 
                    (N577)? 1'b0 : 
                    (N75)? 1'b1 : 
                    (N76)? 1'b1 : 
                    (N77)? 1'b1 : 
                    (N78)? 1'b1 : 
                    (N79)? 1'b0 : 
                    (N80)? 1'b0 : 
                    (N81)? 1'b0 : 
                    (N82)? 1'b0 : 
                    (N83)? 1'b1 : 
                    (N84)? 1'b1 : 
                    (N85)? 1'b1 : 
                    (N648)? 1'b1 : 
                    (N86)? 1'b0 : 
                    (N87)? 1'b0 : 
                    (N88)? 1'b0 : 
                    (N678)? 1'b0 : 
                    (N89)? 1'b1 : 
                    (N90)? 1'b1 : 
                    (N91)? 1'b1 : 
                    (N92)? 1'b0 : 
                    (N93)? 1'b0 : 
                    (N94)? 1'b0 : 
                    (N95)? 1'b0 : 
                    (N96)? 1'b1 : 
                    (N97)? 1'b1 : 
                    (N98)? 1'b1 : 
                    (N740)? 1'b1 : 
                    (N99)? 1'b0 : 
                    (N100)? 1'b0 : 
                    (N101)? 1'b0 : 
                    (N102)? 1'b0 : 
                    (N792)? 1'b1 : 
                    (N103)? 1'b1 : 
                    (N104)? 1'b1 : 
                    (N105)? 1'b0 : 
                    (N106)? 1'b0 : 
                    (N107)? 1'b0 : 
                    (N108)? 1'b0 : 
                    (N109)? 1'b1 : 
                    (N110)? 1'b1 : 
                    (N111)? 1'b1 : 
                    (N848)? 1'b1 : 
                    (N112)? 1'b0 : 
                    (N113)? 1'b0 : 
                    (N114)? 1'b0 : 
                    (N115)? 1'b0 : 
                    (N116)? 1'b1 : 
                    (N898)? 1'b1 : 
                    (N117)? 1'b1 : 
                    (N118)? 1'b0 : 
                    (N119)? 1'b0 : 
                    (N120)? 1'b0 : 
                    (N121)? 1'b0 : 
                    (N122)? 1'b1 : 
                    (N123)? 1'b1 : 
                    (N124)? 1'b1 : 
                    (N948)? 1'b1 : 
                    (N125)? 1'b0 : 
                    (N126)? 1'b0 : 
                    (N127)? 1'b0 : 
                    (N128)? 1'b0 : 
                    (N129)? 1'b1 : 
                    (N130)? 1'b1 : 
                    (N1009)? 1'b1 : 
                    (N131)? 1'b0 : 
                    (N132)? 1'b0 : 
                    (N133)? 1'b0 : 
                    (N134)? 1'b0 : 
                    (N135)? 1'b1 : 
                    (N136)? 1'b1 : 
                    (N137)? 1'b1 : 
                    (N1054)? 1'b1 : 
                    (N138)? 1'b0 : 
                    (N139)? 1'b0 : 
                    (N140)? 1'b0 : 
                    (N141)? 1'b0 : 
                    (N142)? 1'b1 : 
                    (N143)? 1'b1 : 
                    (N144)? 1'b1 : 
                    (N1109)? 1'b1 : 
                    (N145)? 1'b0 : 
                    (N146)? 1'b0 : 
                    (N147)? 1'b0 : 
                    (N148)? 1'b1 : 
                    (N149)? 1'b1 : 
                    (N150)? 1'b1 : 
                    (N1147)? 1'b1 : 
                    (N151)? 1'b0 : 
                    (N152)? 1'b0 : 
                    (N153)? 1'b0 : 
                    (N154)? 1'b0 : 
                    (N155)? 1'b1 : 
                    (N156)? 1'b1 : 
                    (N157)? 1'b1 : 
                    (N158)? 1'b1 : 
                    (N1224)? 1'b0 : 
                    (N159)? 1'b0 : 
                    (N160)? 1'b0 : 
                    (N161)? 1'b1 : 
                    (N162)? 1'b1 : 
                    (N163)? 1'b1 : 
                    (N1256)? 1'b1 : 
                    (N164)? 1'b0 : 
                    (N165)? 1'b0 : 
                    (N166)? 1'b0 : 
                    (N167)? 1'b0 : 
                    (N168)? 1'b1 : 
                    (N169)? 1'b1 : 
                    (N170)? 1'b1 : 
                    (N171)? 1'b1 : 
                    (N172)? 1'b0 : 
                    (N1330)? 1'b0 : 
                    (N173)? 1'b0 : 
                    (N174)? 1'b1 : 
                    (N175)? 1'b1 : 
                    (N176)? 1'b1 : 
                    (N1356)? 1'b1 : 
                    (N177)? 1'b0 : 
                    (N178)? 1'b0 : 
                    (N179)? 1'b0 : 
                    (N180)? 1'b0 : 
                    (N181)? 1'b1 : 
                    (N182)? 1'b1 : 
                    (N183)? 1'b1 : 
                    (N184)? 1'b1 : 
                    (N185)? 1'b0 : 
                    (N186)? 1'b0 : 
                    (N1446)? 1'b0 : 
                    (N187)? 1'b1 : 
                    (N188)? 1'b1 : 
                    (N189)? 1'b1 : 
                    (N1468)? 1'b1 : 
                    (N190)? 1'b0 : 
                    (N191)? 1'b0 : 
                    (N192)? 1'b0 : 
                    (N193)? 1'b0 : 
                    (N194)? 1'b1 : 
                    (N195)? 1'b1 : 
                    (N196)? 1'b1 : 
                    (N197)? 1'b1 : 
                    (N198)? 1'b0 : 
                    (N199)? 1'b0 : 
                    (N200)? 1'b0 : 
                    (N1547)? 1'b0 : 
                    (N201)? 1'b1 : 
                    (N202)? 1'b1 : 
                    (N1563)? 1'b1 : 
                    (N203)? 1'b0 : 
                    (N204)? 1'b0 : 
                    (N205)? 1'b0 : 
                    (N206)? 1'b0 : 
                    (N207)? 1'b1 : 
                    (N208)? 1'b1 : 
                    (N209)? 1'b1 : 
                    (N210)? 1'b1 : 
                    (N211)? 1'b0 : 
                    (N212)? 1'b0 : 
                    (N213)? 1'b0 : 
                    (N214)? 1'b0 : 
                    (N1665)? 1'b1 : 
                    (N215)? 1'b1 : 
                    (N1675)? 1'b1 : 
                    (N216)? 1'b0 : 
                    (N217)? 1'b0 : 
                    (N218)? 1'b0 : 
                    (N219)? 1'b0 : 
                    (N220)? 1'b1 : 
                    (N221)? 1'b1 : 
                    (N222)? 1'b1 : 
                    (N223)? 1'b1 : 
                    (N224)? 1'b0 : 
                    (N225)? 1'b0 : 
                    (N226)? 1'b0 : 
                    (N227)? 1'b0 : 
                    (N228)? 1'b1 : 
                    (N1763)? 1'b1 : 
                    (N1768)? 1'b1 : 
                    (N229)? 1'b0 : 
                    (N230)? 1'b0 : 
                    (N231)? 1'b0 : 
                    (N232)? 1'b0 : 
                    (N233)? 1'b1 : 
                    (N234)? 1'b1 : 
                    (N235)? 1'b1 : 
                    (N236)? 1'b1 : 
                    (N237)? 1'b0 : 
                    (N238)? 1'b0 : 
                    (N239)? 1'b0 : 
                    (N240)? 1'b0 : 
                    (N241)? 1'b1 : 
                    (N242)? 1'b1 : 
                    (N1874)? 1'b1 : 
                    (N243)? 1'b0 : 
                    (N244)? 1'b0 : 
                    (N245)? 1'b0 : 
                    (N246)? 1'b0 : 
                    (N247)? 1'b1 : 
                    (N248)? 1'b1 : 
                    (N249)? 1'b1 : 
                    (N250)? 1'b1 : 
                    (N251)? 1'b0 : 
                    (N252)? 1'b0 : 
                    (N253)? 1'b0 : 
                    (N254)? 1'b0 : 
                    (N255)? 1'b1 : 
                    (N256)? 1'b1 : 
                    (N257)? 1'b1 : 
                    (N1957)? 1'b1 : 1'b0;
  assign tag_o[1] = (N32)? 1'b0 : 
                    (N33)? 1'b0 : 
                    (N34)? 1'b1 : 
                    (N35)? 1'b1 : 
                    (N36)? 1'b0 : 
                    (N37)? 1'b0 : 
                    (N38)? 1'b1 : 
                    (N39)? 1'b1 : 
                    (N40)? 1'b0 : 
                    (N41)? 1'b0 : 
                    (N42)? 1'b1 : 
                    (N43)? 1'b1 : 
                    (N44)? 1'b0 : 
                    (N45)? 1'b0 : 
                    (N46)? 1'b1 : 
                    (N371)? 1'b1 : 
                    (N382)? 1'b0 : 
                    (N47)? 1'b1 : 
                    (N48)? 1'b1 : 
                    (N49)? 1'b0 : 
                    (N50)? 1'b0 : 
                    (N51)? 1'b1 : 
                    (N52)? 1'b1 : 
                    (N53)? 1'b0 : 
                    (N54)? 1'b0 : 
                    (N55)? 1'b1 : 
                    (N56)? 1'b1 : 
                    (N57)? 1'b0 : 
                    (N58)? 1'b0 : 
                    (N59)? 1'b1 : 
                    (N462)? 1'b1 : 
                    (N60)? 1'b0 : 
                    (N479)? 1'b0 : 
                    (N61)? 1'b1 : 
                    (N62)? 1'b0 : 
                    (N63)? 1'b0 : 
                    (N64)? 1'b1 : 
                    (N65)? 1'b1 : 
                    (N66)? 1'b0 : 
                    (N67)? 1'b0 : 
                    (N68)? 1'b1 : 
                    (N69)? 1'b1 : 
                    (N70)? 1'b0 : 
                    (N71)? 1'b0 : 
                    (N72)? 1'b1 : 
                    (N552)? 1'b1 : 
                    (N73)? 1'b0 : 
                    (N74)? 1'b0 : 
                    (N577)? 1'b1 : 
                    (N75)? 1'b0 : 
                    (N76)? 1'b0 : 
                    (N77)? 1'b1 : 
                    (N78)? 1'b1 : 
                    (N79)? 1'b0 : 
                    (N80)? 1'b0 : 
                    (N81)? 1'b1 : 
                    (N82)? 1'b1 : 
                    (N83)? 1'b0 : 
                    (N84)? 1'b0 : 
                    (N85)? 1'b1 : 
                    (N648)? 1'b1 : 
                    (N86)? 1'b0 : 
                    (N87)? 1'b0 : 
                    (N88)? 1'b1 : 
                    (N678)? 1'b1 : 
                    (N89)? 1'b0 : 
                    (N90)? 1'b1 : 
                    (N91)? 1'b1 : 
                    (N92)? 1'b0 : 
                    (N93)? 1'b0 : 
                    (N94)? 1'b1 : 
                    (N95)? 1'b1 : 
                    (N96)? 1'b0 : 
                    (N97)? 1'b0 : 
                    (N98)? 1'b1 : 
                    (N740)? 1'b1 : 
                    (N99)? 1'b0 : 
                    (N100)? 1'b0 : 
                    (N101)? 1'b1 : 
                    (N102)? 1'b1 : 
                    (N792)? 1'b0 : 
                    (N103)? 1'b1 : 
                    (N104)? 1'b1 : 
                    (N105)? 1'b0 : 
                    (N106)? 1'b0 : 
                    (N107)? 1'b1 : 
                    (N108)? 1'b1 : 
                    (N109)? 1'b0 : 
                    (N110)? 1'b0 : 
                    (N111)? 1'b1 : 
                    (N848)? 1'b1 : 
                    (N112)? 1'b0 : 
                    (N113)? 1'b0 : 
                    (N114)? 1'b1 : 
                    (N115)? 1'b1 : 
                    (N116)? 1'b0 : 
                    (N898)? 1'b0 : 
                    (N117)? 1'b1 : 
                    (N118)? 1'b0 : 
                    (N119)? 1'b0 : 
                    (N120)? 1'b1 : 
                    (N121)? 1'b1 : 
                    (N122)? 1'b0 : 
                    (N123)? 1'b0 : 
                    (N124)? 1'b1 : 
                    (N948)? 1'b1 : 
                    (N125)? 1'b0 : 
                    (N126)? 1'b0 : 
                    (N127)? 1'b1 : 
                    (N128)? 1'b1 : 
                    (N129)? 1'b0 : 
                    (N130)? 1'b0 : 
                    (N1009)? 1'b1 : 
                    (N131)? 1'b0 : 
                    (N132)? 1'b0 : 
                    (N133)? 1'b1 : 
                    (N134)? 1'b1 : 
                    (N135)? 1'b0 : 
                    (N136)? 1'b0 : 
                    (N137)? 1'b1 : 
                    (N1054)? 1'b1 : 
                    (N138)? 1'b0 : 
                    (N139)? 1'b0 : 
                    (N140)? 1'b1 : 
                    (N141)? 1'b1 : 
                    (N142)? 1'b0 : 
                    (N143)? 1'b0 : 
                    (N144)? 1'b1 : 
                    (N1109)? 1'b1 : 
                    (N145)? 1'b0 : 
                    (N146)? 1'b1 : 
                    (N147)? 1'b1 : 
                    (N148)? 1'b0 : 
                    (N149)? 1'b0 : 
                    (N150)? 1'b1 : 
                    (N1147)? 1'b1 : 
                    (N151)? 1'b0 : 
                    (N152)? 1'b0 : 
                    (N153)? 1'b1 : 
                    (N154)? 1'b1 : 
                    (N155)? 1'b0 : 
                    (N156)? 1'b0 : 
                    (N157)? 1'b1 : 
                    (N158)? 1'b1 : 
                    (N1224)? 1'b0 : 
                    (N159)? 1'b1 : 
                    (N160)? 1'b1 : 
                    (N161)? 1'b0 : 
                    (N162)? 1'b0 : 
                    (N163)? 1'b1 : 
                    (N1256)? 1'b1 : 
                    (N164)? 1'b0 : 
                    (N165)? 1'b0 : 
                    (N166)? 1'b1 : 
                    (N167)? 1'b1 : 
                    (N168)? 1'b0 : 
                    (N169)? 1'b0 : 
                    (N170)? 1'b1 : 
                    (N171)? 1'b1 : 
                    (N172)? 1'b0 : 
                    (N1330)? 1'b0 : 
                    (N173)? 1'b1 : 
                    (N174)? 1'b0 : 
                    (N175)? 1'b0 : 
                    (N176)? 1'b1 : 
                    (N1356)? 1'b1 : 
                    (N177)? 1'b0 : 
                    (N178)? 1'b0 : 
                    (N179)? 1'b1 : 
                    (N180)? 1'b1 : 
                    (N181)? 1'b0 : 
                    (N182)? 1'b0 : 
                    (N183)? 1'b1 : 
                    (N184)? 1'b1 : 
                    (N185)? 1'b0 : 
                    (N186)? 1'b0 : 
                    (N1446)? 1'b1 : 
                    (N187)? 1'b0 : 
                    (N188)? 1'b0 : 
                    (N189)? 1'b1 : 
                    (N1468)? 1'b1 : 
                    (N190)? 1'b0 : 
                    (N191)? 1'b0 : 
                    (N192)? 1'b1 : 
                    (N193)? 1'b1 : 
                    (N194)? 1'b0 : 
                    (N195)? 1'b0 : 
                    (N196)? 1'b1 : 
                    (N197)? 1'b1 : 
                    (N198)? 1'b0 : 
                    (N199)? 1'b0 : 
                    (N200)? 1'b1 : 
                    (N1547)? 1'b1 : 
                    (N201)? 1'b0 : 
                    (N202)? 1'b1 : 
                    (N1563)? 1'b1 : 
                    (N203)? 1'b0 : 
                    (N204)? 1'b0 : 
                    (N205)? 1'b1 : 
                    (N206)? 1'b1 : 
                    (N207)? 1'b0 : 
                    (N208)? 1'b0 : 
                    (N209)? 1'b1 : 
                    (N210)? 1'b1 : 
                    (N211)? 1'b0 : 
                    (N212)? 1'b0 : 
                    (N213)? 1'b1 : 
                    (N214)? 1'b1 : 
                    (N1665)? 1'b0 : 
                    (N215)? 1'b1 : 
                    (N1675)? 1'b1 : 
                    (N216)? 1'b0 : 
                    (N217)? 1'b0 : 
                    (N218)? 1'b1 : 
                    (N219)? 1'b1 : 
                    (N220)? 1'b0 : 
                    (N221)? 1'b0 : 
                    (N222)? 1'b1 : 
                    (N223)? 1'b1 : 
                    (N224)? 1'b0 : 
                    (N225)? 1'b0 : 
                    (N226)? 1'b1 : 
                    (N227)? 1'b1 : 
                    (N228)? 1'b0 : 
                    (N1763)? 1'b0 : 
                    (N1768)? 1'b1 : 
                    (N229)? 1'b0 : 
                    (N230)? 1'b0 : 
                    (N231)? 1'b1 : 
                    (N232)? 1'b1 : 
                    (N233)? 1'b0 : 
                    (N234)? 1'b0 : 
                    (N235)? 1'b1 : 
                    (N236)? 1'b1 : 
                    (N237)? 1'b0 : 
                    (N238)? 1'b0 : 
                    (N239)? 1'b1 : 
                    (N240)? 1'b1 : 
                    (N241)? 1'b0 : 
                    (N242)? 1'b0 : 
                    (N1874)? 1'b1 : 
                    (N243)? 1'b0 : 
                    (N244)? 1'b0 : 
                    (N245)? 1'b1 : 
                    (N246)? 1'b1 : 
                    (N247)? 1'b0 : 
                    (N248)? 1'b0 : 
                    (N249)? 1'b1 : 
                    (N250)? 1'b1 : 
                    (N251)? 1'b0 : 
                    (N252)? 1'b0 : 
                    (N253)? 1'b1 : 
                    (N254)? 1'b1 : 
                    (N255)? 1'b0 : 
                    (N256)? 1'b0 : 
                    (N257)? 1'b1 : 
                    (N1957)? 1'b1 : 1'b0;
  assign tag_o[0] = (N32)? 1'b0 : 
                    (N33)? 1'b1 : 
                    (N34)? 1'b0 : 
                    (N35)? 1'b1 : 
                    (N36)? 1'b0 : 
                    (N37)? 1'b1 : 
                    (N38)? 1'b0 : 
                    (N39)? 1'b1 : 
                    (N40)? 1'b0 : 
                    (N41)? 1'b1 : 
                    (N42)? 1'b0 : 
                    (N43)? 1'b1 : 
                    (N44)? 1'b0 : 
                    (N45)? 1'b1 : 
                    (N46)? 1'b0 : 
                    (N371)? 1'b1 : 
                    (N382)? 1'b0 : 
                    (N47)? 1'b0 : 
                    (N48)? 1'b1 : 
                    (N49)? 1'b0 : 
                    (N50)? 1'b1 : 
                    (N51)? 1'b0 : 
                    (N52)? 1'b1 : 
                    (N53)? 1'b0 : 
                    (N54)? 1'b1 : 
                    (N55)? 1'b0 : 
                    (N56)? 1'b1 : 
                    (N57)? 1'b0 : 
                    (N58)? 1'b1 : 
                    (N59)? 1'b0 : 
                    (N462)? 1'b1 : 
                    (N60)? 1'b0 : 
                    (N479)? 1'b1 : 
                    (N61)? 1'b1 : 
                    (N62)? 1'b0 : 
                    (N63)? 1'b1 : 
                    (N64)? 1'b0 : 
                    (N65)? 1'b1 : 
                    (N66)? 1'b0 : 
                    (N67)? 1'b1 : 
                    (N68)? 1'b0 : 
                    (N69)? 1'b1 : 
                    (N70)? 1'b0 : 
                    (N71)? 1'b1 : 
                    (N72)? 1'b0 : 
                    (N552)? 1'b1 : 
                    (N73)? 1'b0 : 
                    (N74)? 1'b1 : 
                    (N577)? 1'b0 : 
                    (N75)? 1'b0 : 
                    (N76)? 1'b1 : 
                    (N77)? 1'b0 : 
                    (N78)? 1'b1 : 
                    (N79)? 1'b0 : 
                    (N80)? 1'b1 : 
                    (N81)? 1'b0 : 
                    (N82)? 1'b1 : 
                    (N83)? 1'b0 : 
                    (N84)? 1'b1 : 
                    (N85)? 1'b0 : 
                    (N648)? 1'b1 : 
                    (N86)? 1'b0 : 
                    (N87)? 1'b1 : 
                    (N88)? 1'b0 : 
                    (N678)? 1'b1 : 
                    (N89)? 1'b1 : 
                    (N90)? 1'b0 : 
                    (N91)? 1'b1 : 
                    (N92)? 1'b0 : 
                    (N93)? 1'b1 : 
                    (N94)? 1'b0 : 
                    (N95)? 1'b1 : 
                    (N96)? 1'b0 : 
                    (N97)? 1'b1 : 
                    (N98)? 1'b0 : 
                    (N740)? 1'b1 : 
                    (N99)? 1'b0 : 
                    (N100)? 1'b1 : 
                    (N101)? 1'b0 : 
                    (N102)? 1'b1 : 
                    (N792)? 1'b0 : 
                    (N103)? 1'b0 : 
                    (N104)? 1'b1 : 
                    (N105)? 1'b0 : 
                    (N106)? 1'b1 : 
                    (N107)? 1'b0 : 
                    (N108)? 1'b1 : 
                    (N109)? 1'b0 : 
                    (N110)? 1'b1 : 
                    (N111)? 1'b0 : 
                    (N848)? 1'b1 : 
                    (N112)? 1'b0 : 
                    (N113)? 1'b1 : 
                    (N114)? 1'b0 : 
                    (N115)? 1'b1 : 
                    (N116)? 1'b0 : 
                    (N898)? 1'b1 : 
                    (N117)? 1'b1 : 
                    (N118)? 1'b0 : 
                    (N119)? 1'b1 : 
                    (N120)? 1'b0 : 
                    (N121)? 1'b1 : 
                    (N122)? 1'b0 : 
                    (N123)? 1'b1 : 
                    (N124)? 1'b0 : 
                    (N948)? 1'b1 : 
                    (N125)? 1'b0 : 
                    (N126)? 1'b1 : 
                    (N127)? 1'b0 : 
                    (N128)? 1'b1 : 
                    (N129)? 1'b0 : 
                    (N130)? 1'b1 : 
                    (N1009)? 1'b0 : 
                    (N131)? 1'b0 : 
                    (N132)? 1'b1 : 
                    (N133)? 1'b0 : 
                    (N134)? 1'b1 : 
                    (N135)? 1'b0 : 
                    (N136)? 1'b1 : 
                    (N137)? 1'b0 : 
                    (N1054)? 1'b1 : 
                    (N138)? 1'b0 : 
                    (N139)? 1'b1 : 
                    (N140)? 1'b0 : 
                    (N141)? 1'b1 : 
                    (N142)? 1'b0 : 
                    (N143)? 1'b1 : 
                    (N144)? 1'b0 : 
                    (N1109)? 1'b1 : 
                    (N145)? 1'b1 : 
                    (N146)? 1'b0 : 
                    (N147)? 1'b1 : 
                    (N148)? 1'b0 : 
                    (N149)? 1'b1 : 
                    (N150)? 1'b0 : 
                    (N1147)? 1'b1 : 
                    (N151)? 1'b0 : 
                    (N152)? 1'b1 : 
                    (N153)? 1'b0 : 
                    (N154)? 1'b1 : 
                    (N155)? 1'b0 : 
                    (N156)? 1'b1 : 
                    (N157)? 1'b0 : 
                    (N158)? 1'b1 : 
                    (N1224)? 1'b0 : 
                    (N159)? 1'b0 : 
                    (N160)? 1'b1 : 
                    (N161)? 1'b0 : 
                    (N162)? 1'b1 : 
                    (N163)? 1'b0 : 
                    (N1256)? 1'b1 : 
                    (N164)? 1'b0 : 
                    (N165)? 1'b1 : 
                    (N166)? 1'b0 : 
                    (N167)? 1'b1 : 
                    (N168)? 1'b0 : 
                    (N169)? 1'b1 : 
                    (N170)? 1'b0 : 
                    (N171)? 1'b1 : 
                    (N172)? 1'b0 : 
                    (N1330)? 1'b1 : 
                    (N173)? 1'b1 : 
                    (N174)? 1'b0 : 
                    (N175)? 1'b1 : 
                    (N176)? 1'b0 : 
                    (N1356)? 1'b1 : 
                    (N177)? 1'b0 : 
                    (N178)? 1'b1 : 
                    (N179)? 1'b0 : 
                    (N180)? 1'b1 : 
                    (N181)? 1'b0 : 
                    (N182)? 1'b1 : 
                    (N183)? 1'b0 : 
                    (N184)? 1'b1 : 
                    (N185)? 1'b0 : 
                    (N186)? 1'b1 : 
                    (N1446)? 1'b0 : 
                    (N187)? 1'b0 : 
                    (N188)? 1'b1 : 
                    (N189)? 1'b0 : 
                    (N1468)? 1'b1 : 
                    (N190)? 1'b0 : 
                    (N191)? 1'b1 : 
                    (N192)? 1'b0 : 
                    (N193)? 1'b1 : 
                    (N194)? 1'b0 : 
                    (N195)? 1'b1 : 
                    (N196)? 1'b0 : 
                    (N197)? 1'b1 : 
                    (N198)? 1'b0 : 
                    (N199)? 1'b1 : 
                    (N200)? 1'b0 : 
                    (N1547)? 1'b1 : 
                    (N201)? 1'b1 : 
                    (N202)? 1'b0 : 
                    (N1563)? 1'b1 : 
                    (N203)? 1'b0 : 
                    (N204)? 1'b1 : 
                    (N205)? 1'b0 : 
                    (N206)? 1'b1 : 
                    (N207)? 1'b0 : 
                    (N208)? 1'b1 : 
                    (N209)? 1'b0 : 
                    (N210)? 1'b1 : 
                    (N211)? 1'b0 : 
                    (N212)? 1'b1 : 
                    (N213)? 1'b0 : 
                    (N214)? 1'b1 : 
                    (N1665)? 1'b0 : 
                    (N215)? 1'b0 : 
                    (N1675)? 1'b1 : 
                    (N216)? 1'b0 : 
                    (N217)? 1'b1 : 
                    (N218)? 1'b0 : 
                    (N219)? 1'b1 : 
                    (N220)? 1'b0 : 
                    (N221)? 1'b1 : 
                    (N222)? 1'b0 : 
                    (N223)? 1'b1 : 
                    (N224)? 1'b0 : 
                    (N225)? 1'b1 : 
                    (N226)? 1'b0 : 
                    (N227)? 1'b1 : 
                    (N228)? 1'b0 : 
                    (N1763)? 1'b1 : 
                    (N1768)? 1'b1 : 
                    (N229)? 1'b0 : 
                    (N230)? 1'b1 : 
                    (N231)? 1'b0 : 
                    (N232)? 1'b1 : 
                    (N233)? 1'b0 : 
                    (N234)? 1'b1 : 
                    (N235)? 1'b0 : 
                    (N236)? 1'b1 : 
                    (N237)? 1'b0 : 
                    (N238)? 1'b1 : 
                    (N239)? 1'b0 : 
                    (N240)? 1'b1 : 
                    (N241)? 1'b0 : 
                    (N242)? 1'b1 : 
                    (N1874)? 1'b0 : 
                    (N243)? 1'b0 : 
                    (N244)? 1'b1 : 
                    (N245)? 1'b0 : 
                    (N246)? 1'b1 : 
                    (N247)? 1'b0 : 
                    (N248)? 1'b1 : 
                    (N249)? 1'b0 : 
                    (N250)? 1'b1 : 
                    (N251)? 1'b0 : 
                    (N252)? 1'b1 : 
                    (N253)? 1'b0 : 
                    (N254)? 1'b1 : 
                    (N255)? 1'b0 : 
                    (N256)? 1'b1 : 
                    (N257)? 1'b0 : 
                    (N1957)? 1'b1 : 1'b0;
  assign N258 = ~reqs_i[6];
  assign N259 = ~reqs_i[5];
  assign N260 = ~reqs_i[4];
  assign N270 = ~last_r[3];
  assign N271 = ~last_r[2];
  assign N272 = ~last_r[1];
  assign N273 = ~last_r[0];
  assign N278 = ~reqs_i[1];
  assign N290 = ~reqs_i[3];
  assign N304 = ~reqs_i[2];
  assign N371 = ~N370;
  assign N382 = ~N381;
  assign N462 = ~N461;
  assign N479 = ~N478;
  assign N552 = ~N551;
  assign N560 = ~reqs_i[0];
  assign N577 = ~N576;
  assign N648 = ~N647;
  assign N678 = ~N677;
  assign N740 = ~N739;
  assign N741 = ~reqs_i[15];
  assign N792 = ~N791;
  assign N848 = ~N847;
  assign N898 = ~N897;
  assign N918 = ~reqs_i[7];
  assign N948 = ~N947;
  assign N1009 = ~N1008;
  assign N1029 = ~reqs_i[8];
  assign N1054 = ~N1053;
  assign N1109 = ~N1108;
  assign N1129 = ~reqs_i[9];
  assign N1147 = ~N1146;
  assign N1224 = ~N1223;
  assign N1244 = ~reqs_i[10];
  assign N1256 = ~N1255;
  assign N1330 = ~N1329;
  assign N1356 = ~N1355;
  assign N1357 = ~reqs_i[11];
  assign N1446 = ~N1445;
  assign N1451 = ~reqs_i[12];
  assign N1468 = ~N1467;
  assign N1547 = ~N1546;
  assign N1552 = ~reqs_i[13];
  assign N1563 = ~N1562;
  assign N1564 = ~reqs_i[14];
  assign N1665 = ~N1664;
  assign N1675 = ~N1674;
  assign N1763 = ~N1762;
  assign N1768 = ~N1767;
  assign N1874 = ~N1873;
  assign N1957 = ~N1956;
  assign grants_o[15] = sel_one_hot_o[15] & grants_en_i;
  assign grants_o[14] = sel_one_hot_o[14] & grants_en_i;
  assign grants_o[13] = sel_one_hot_o[13] & grants_en_i;
  assign grants_o[12] = sel_one_hot_o[12] & grants_en_i;
  assign grants_o[11] = sel_one_hot_o[11] & grants_en_i;
  assign grants_o[10] = sel_one_hot_o[10] & grants_en_i;
  assign grants_o[9] = sel_one_hot_o[9] & grants_en_i;
  assign grants_o[8] = sel_one_hot_o[8] & grants_en_i;
  assign grants_o[7] = sel_one_hot_o[7] & grants_en_i;
  assign grants_o[6] = sel_one_hot_o[6] & grants_en_i;
  assign grants_o[5] = sel_one_hot_o[5] & grants_en_i;
  assign grants_o[4] = sel_one_hot_o[4] & grants_en_i;
  assign grants_o[3] = sel_one_hot_o[3] & grants_en_i;
  assign grants_o[2] = sel_one_hot_o[2] & grants_en_i;
  assign grants_o[1] = sel_one_hot_o[1] & grants_en_i;
  assign grants_o[0] = sel_one_hot_o[0] & grants_en_i;
  assign v_o = N2530 | reqs_i[0];
  assign N2530 = N2529 | reqs_i[1];
  assign N2529 = N2528 | reqs_i[2];
  assign N2528 = N2527 | reqs_i[3];
  assign N2527 = N2526 | reqs_i[4];
  assign N2526 = N2525 | reqs_i[5];
  assign N2525 = N2524 | reqs_i[6];
  assign N2524 = N2523 | reqs_i[7];
  assign N2523 = N2522 | reqs_i[8];
  assign N2522 = N2521 | reqs_i[9];
  assign N2521 = N2520 | reqs_i[10];
  assign N2520 = N2519 | reqs_i[11];
  assign N2519 = N2518 | reqs_i[12];
  assign N2518 = N2517 | reqs_i[13];
  assign N2517 = reqs_i[15] | reqs_i[14];

  always @(posedge clk_i) begin
    if(reset_i) begin
      last_r_3_sv2v_reg <= 1'b0;
      last_r_2_sv2v_reg <= 1'b0;
      last_r_1_sv2v_reg <= 1'b0;
      last_r_0_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      last_r_3_sv2v_reg <= tag_o[3];
      last_r_2_sv2v_reg <= tag_o[2];
      last_r_1_sv2v_reg <= tag_o[1];
      last_r_0_sv2v_reg <= tag_o[0];
    end 
  end


endmodule

