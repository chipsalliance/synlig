module top(output int o);
   parameter int unsigned P = 20;
   assign o = P;
endmodule
