module top(output shortint o);
   assign o = 1;
endmodule
