
module dut(input logic clk);

localparam int GW_CONFIG2[2:0] = '{default:0} ;

endmodule
