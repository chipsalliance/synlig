module top(output logic a);
   initial begin
      a  = 1; 
      a ^= 0;
   end
endmodule
