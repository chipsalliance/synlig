

module top
(
  i,
  sel_oi_one_hot_i,
  o
);

  input [255:0] i;
  input [255:0] sel_oi_one_hot_i;
  output [255:0] o;

  bsg_crossbar_o_by_i
  wrapper
  (
    .i(i),
    .sel_oi_one_hot_i(sel_oi_one_hot_i),
    .o(o)
  );


endmodule



module bsg_mux_one_hot_width_p16_els_p16
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [255:0] data_i;
  input [15:0] sel_one_hot_i;
  output [15:0] data_o;
  wire [15:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223;
  wire [255:0] data_masked;
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[1];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[1];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[1];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[1];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[1];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[1];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[1];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[1];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[1];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[1];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[1];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[1];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[1];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[1];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[1];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[1];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[2];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[2];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[2];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[2];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[2];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[2];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[2];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[2];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[2];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[2];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[2];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[2];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[2];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[2];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[2];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[2];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[3];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[3];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[3];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[3];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[3];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[3];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[3];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[3];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[3];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[3];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[3];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[3];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[3];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[3];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[3];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[3];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[4];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[4];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[4];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[4];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[4];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[4];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[4];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[4];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[4];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[4];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[4];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[4];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[4];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[4];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[4];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[4];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[5];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[5];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[5];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[5];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[5];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[5];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[5];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[5];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[5];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[5];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[5];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[5];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[5];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[5];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[5];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[5];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[6];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[6];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[6];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[6];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[6];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[6];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[6];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[6];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[6];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[6];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[6];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[6];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[6];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[6];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[6];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[6];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[7];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[7];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[7];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[7];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[7];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[7];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[7];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[7];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[7];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[7];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[7];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[7];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[7];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[7];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[7];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[7];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[8];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[8];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[8];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[8];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[8];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[8];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[8];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[8];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[8];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[8];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[8];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[8];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[8];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[8];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[8];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[8];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[9];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[9];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[9];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[9];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[9];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[9];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[9];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[9];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[9];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[9];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[9];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[9];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[9];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[9];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[9];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[9];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[10];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[10];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[10];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[10];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[10];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[10];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[10];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[10];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[10];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[10];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[10];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[10];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[10];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[10];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[10];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[10];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[11];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[11];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[11];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[11];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[11];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[11];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[11];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[11];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[11];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[11];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[11];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[11];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[11];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[11];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[11];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[11];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[12];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[12];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[12];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[12];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[12];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[12];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[12];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[12];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[12];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[12];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[12];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[12];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[12];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[12];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[12];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[12];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[13];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[13];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[13];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[13];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[13];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[13];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[13];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[13];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[13];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[13];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[13];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[13];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[13];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[13];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[13];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[13];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[14];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[14];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[14];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[14];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[14];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[14];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[14];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[14];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[14];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[14];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[14];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[14];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[14];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[14];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[14];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[14];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[15];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[15];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[15];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[15];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[15];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[15];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[15];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[15];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[15];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[15];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[15];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[15];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[15];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[15];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[15];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[15];
  assign data_o[0] = N13 | data_masked[0];
  assign N13 = N12 | data_masked[16];
  assign N12 = N11 | data_masked[32];
  assign N11 = N10 | data_masked[48];
  assign N10 = N9 | data_masked[64];
  assign N9 = N8 | data_masked[80];
  assign N8 = N7 | data_masked[96];
  assign N7 = N6 | data_masked[112];
  assign N6 = N5 | data_masked[128];
  assign N5 = N4 | data_masked[144];
  assign N4 = N3 | data_masked[160];
  assign N3 = N2 | data_masked[176];
  assign N2 = N1 | data_masked[192];
  assign N1 = N0 | data_masked[208];
  assign N0 = data_masked[240] | data_masked[224];
  assign data_o[1] = N27 | data_masked[1];
  assign N27 = N26 | data_masked[17];
  assign N26 = N25 | data_masked[33];
  assign N25 = N24 | data_masked[49];
  assign N24 = N23 | data_masked[65];
  assign N23 = N22 | data_masked[81];
  assign N22 = N21 | data_masked[97];
  assign N21 = N20 | data_masked[113];
  assign N20 = N19 | data_masked[129];
  assign N19 = N18 | data_masked[145];
  assign N18 = N17 | data_masked[161];
  assign N17 = N16 | data_masked[177];
  assign N16 = N15 | data_masked[193];
  assign N15 = N14 | data_masked[209];
  assign N14 = data_masked[241] | data_masked[225];
  assign data_o[2] = N41 | data_masked[2];
  assign N41 = N40 | data_masked[18];
  assign N40 = N39 | data_masked[34];
  assign N39 = N38 | data_masked[50];
  assign N38 = N37 | data_masked[66];
  assign N37 = N36 | data_masked[82];
  assign N36 = N35 | data_masked[98];
  assign N35 = N34 | data_masked[114];
  assign N34 = N33 | data_masked[130];
  assign N33 = N32 | data_masked[146];
  assign N32 = N31 | data_masked[162];
  assign N31 = N30 | data_masked[178];
  assign N30 = N29 | data_masked[194];
  assign N29 = N28 | data_masked[210];
  assign N28 = data_masked[242] | data_masked[226];
  assign data_o[3] = N55 | data_masked[3];
  assign N55 = N54 | data_masked[19];
  assign N54 = N53 | data_masked[35];
  assign N53 = N52 | data_masked[51];
  assign N52 = N51 | data_masked[67];
  assign N51 = N50 | data_masked[83];
  assign N50 = N49 | data_masked[99];
  assign N49 = N48 | data_masked[115];
  assign N48 = N47 | data_masked[131];
  assign N47 = N46 | data_masked[147];
  assign N46 = N45 | data_masked[163];
  assign N45 = N44 | data_masked[179];
  assign N44 = N43 | data_masked[195];
  assign N43 = N42 | data_masked[211];
  assign N42 = data_masked[243] | data_masked[227];
  assign data_o[4] = N69 | data_masked[4];
  assign N69 = N68 | data_masked[20];
  assign N68 = N67 | data_masked[36];
  assign N67 = N66 | data_masked[52];
  assign N66 = N65 | data_masked[68];
  assign N65 = N64 | data_masked[84];
  assign N64 = N63 | data_masked[100];
  assign N63 = N62 | data_masked[116];
  assign N62 = N61 | data_masked[132];
  assign N61 = N60 | data_masked[148];
  assign N60 = N59 | data_masked[164];
  assign N59 = N58 | data_masked[180];
  assign N58 = N57 | data_masked[196];
  assign N57 = N56 | data_masked[212];
  assign N56 = data_masked[244] | data_masked[228];
  assign data_o[5] = N83 | data_masked[5];
  assign N83 = N82 | data_masked[21];
  assign N82 = N81 | data_masked[37];
  assign N81 = N80 | data_masked[53];
  assign N80 = N79 | data_masked[69];
  assign N79 = N78 | data_masked[85];
  assign N78 = N77 | data_masked[101];
  assign N77 = N76 | data_masked[117];
  assign N76 = N75 | data_masked[133];
  assign N75 = N74 | data_masked[149];
  assign N74 = N73 | data_masked[165];
  assign N73 = N72 | data_masked[181];
  assign N72 = N71 | data_masked[197];
  assign N71 = N70 | data_masked[213];
  assign N70 = data_masked[245] | data_masked[229];
  assign data_o[6] = N97 | data_masked[6];
  assign N97 = N96 | data_masked[22];
  assign N96 = N95 | data_masked[38];
  assign N95 = N94 | data_masked[54];
  assign N94 = N93 | data_masked[70];
  assign N93 = N92 | data_masked[86];
  assign N92 = N91 | data_masked[102];
  assign N91 = N90 | data_masked[118];
  assign N90 = N89 | data_masked[134];
  assign N89 = N88 | data_masked[150];
  assign N88 = N87 | data_masked[166];
  assign N87 = N86 | data_masked[182];
  assign N86 = N85 | data_masked[198];
  assign N85 = N84 | data_masked[214];
  assign N84 = data_masked[246] | data_masked[230];
  assign data_o[7] = N111 | data_masked[7];
  assign N111 = N110 | data_masked[23];
  assign N110 = N109 | data_masked[39];
  assign N109 = N108 | data_masked[55];
  assign N108 = N107 | data_masked[71];
  assign N107 = N106 | data_masked[87];
  assign N106 = N105 | data_masked[103];
  assign N105 = N104 | data_masked[119];
  assign N104 = N103 | data_masked[135];
  assign N103 = N102 | data_masked[151];
  assign N102 = N101 | data_masked[167];
  assign N101 = N100 | data_masked[183];
  assign N100 = N99 | data_masked[199];
  assign N99 = N98 | data_masked[215];
  assign N98 = data_masked[247] | data_masked[231];
  assign data_o[8] = N125 | data_masked[8];
  assign N125 = N124 | data_masked[24];
  assign N124 = N123 | data_masked[40];
  assign N123 = N122 | data_masked[56];
  assign N122 = N121 | data_masked[72];
  assign N121 = N120 | data_masked[88];
  assign N120 = N119 | data_masked[104];
  assign N119 = N118 | data_masked[120];
  assign N118 = N117 | data_masked[136];
  assign N117 = N116 | data_masked[152];
  assign N116 = N115 | data_masked[168];
  assign N115 = N114 | data_masked[184];
  assign N114 = N113 | data_masked[200];
  assign N113 = N112 | data_masked[216];
  assign N112 = data_masked[248] | data_masked[232];
  assign data_o[9] = N139 | data_masked[9];
  assign N139 = N138 | data_masked[25];
  assign N138 = N137 | data_masked[41];
  assign N137 = N136 | data_masked[57];
  assign N136 = N135 | data_masked[73];
  assign N135 = N134 | data_masked[89];
  assign N134 = N133 | data_masked[105];
  assign N133 = N132 | data_masked[121];
  assign N132 = N131 | data_masked[137];
  assign N131 = N130 | data_masked[153];
  assign N130 = N129 | data_masked[169];
  assign N129 = N128 | data_masked[185];
  assign N128 = N127 | data_masked[201];
  assign N127 = N126 | data_masked[217];
  assign N126 = data_masked[249] | data_masked[233];
  assign data_o[10] = N153 | data_masked[10];
  assign N153 = N152 | data_masked[26];
  assign N152 = N151 | data_masked[42];
  assign N151 = N150 | data_masked[58];
  assign N150 = N149 | data_masked[74];
  assign N149 = N148 | data_masked[90];
  assign N148 = N147 | data_masked[106];
  assign N147 = N146 | data_masked[122];
  assign N146 = N145 | data_masked[138];
  assign N145 = N144 | data_masked[154];
  assign N144 = N143 | data_masked[170];
  assign N143 = N142 | data_masked[186];
  assign N142 = N141 | data_masked[202];
  assign N141 = N140 | data_masked[218];
  assign N140 = data_masked[250] | data_masked[234];
  assign data_o[11] = N167 | data_masked[11];
  assign N167 = N166 | data_masked[27];
  assign N166 = N165 | data_masked[43];
  assign N165 = N164 | data_masked[59];
  assign N164 = N163 | data_masked[75];
  assign N163 = N162 | data_masked[91];
  assign N162 = N161 | data_masked[107];
  assign N161 = N160 | data_masked[123];
  assign N160 = N159 | data_masked[139];
  assign N159 = N158 | data_masked[155];
  assign N158 = N157 | data_masked[171];
  assign N157 = N156 | data_masked[187];
  assign N156 = N155 | data_masked[203];
  assign N155 = N154 | data_masked[219];
  assign N154 = data_masked[251] | data_masked[235];
  assign data_o[12] = N181 | data_masked[12];
  assign N181 = N180 | data_masked[28];
  assign N180 = N179 | data_masked[44];
  assign N179 = N178 | data_masked[60];
  assign N178 = N177 | data_masked[76];
  assign N177 = N176 | data_masked[92];
  assign N176 = N175 | data_masked[108];
  assign N175 = N174 | data_masked[124];
  assign N174 = N173 | data_masked[140];
  assign N173 = N172 | data_masked[156];
  assign N172 = N171 | data_masked[172];
  assign N171 = N170 | data_masked[188];
  assign N170 = N169 | data_masked[204];
  assign N169 = N168 | data_masked[220];
  assign N168 = data_masked[252] | data_masked[236];
  assign data_o[13] = N195 | data_masked[13];
  assign N195 = N194 | data_masked[29];
  assign N194 = N193 | data_masked[45];
  assign N193 = N192 | data_masked[61];
  assign N192 = N191 | data_masked[77];
  assign N191 = N190 | data_masked[93];
  assign N190 = N189 | data_masked[109];
  assign N189 = N188 | data_masked[125];
  assign N188 = N187 | data_masked[141];
  assign N187 = N186 | data_masked[157];
  assign N186 = N185 | data_masked[173];
  assign N185 = N184 | data_masked[189];
  assign N184 = N183 | data_masked[205];
  assign N183 = N182 | data_masked[221];
  assign N182 = data_masked[253] | data_masked[237];
  assign data_o[14] = N209 | data_masked[14];
  assign N209 = N208 | data_masked[30];
  assign N208 = N207 | data_masked[46];
  assign N207 = N206 | data_masked[62];
  assign N206 = N205 | data_masked[78];
  assign N205 = N204 | data_masked[94];
  assign N204 = N203 | data_masked[110];
  assign N203 = N202 | data_masked[126];
  assign N202 = N201 | data_masked[142];
  assign N201 = N200 | data_masked[158];
  assign N200 = N199 | data_masked[174];
  assign N199 = N198 | data_masked[190];
  assign N198 = N197 | data_masked[206];
  assign N197 = N196 | data_masked[222];
  assign N196 = data_masked[254] | data_masked[238];
  assign data_o[15] = N223 | data_masked[15];
  assign N223 = N222 | data_masked[31];
  assign N222 = N221 | data_masked[47];
  assign N221 = N220 | data_masked[63];
  assign N220 = N219 | data_masked[79];
  assign N219 = N218 | data_masked[95];
  assign N218 = N217 | data_masked[111];
  assign N217 = N216 | data_masked[127];
  assign N216 = N215 | data_masked[143];
  assign N215 = N214 | data_masked[159];
  assign N214 = N213 | data_masked[175];
  assign N213 = N212 | data_masked[191];
  assign N212 = N211 | data_masked[207];
  assign N211 = N210 | data_masked[223];
  assign N210 = data_masked[255] | data_masked[239];

endmodule



module bsg_crossbar_o_by_i
(
  i,
  sel_oi_one_hot_i,
  o
);

  input [255:0] i;
  input [255:0] sel_oi_one_hot_i;
  output [255:0] o;
  wire [255:0] o;

  bsg_mux_one_hot_width_p16_els_p16
  \l_0_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[15:0]),
    .data_o(o[15:0])
  );


  bsg_mux_one_hot_width_p16_els_p16
  \l_1_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[31:16]),
    .data_o(o[31:16])
  );


  bsg_mux_one_hot_width_p16_els_p16
  \l_2_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[47:32]),
    .data_o(o[47:32])
  );


  bsg_mux_one_hot_width_p16_els_p16
  \l_3_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[63:48]),
    .data_o(o[63:48])
  );


  bsg_mux_one_hot_width_p16_els_p16
  \l_4_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[79:64]),
    .data_o(o[79:64])
  );


  bsg_mux_one_hot_width_p16_els_p16
  \l_5_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[95:80]),
    .data_o(o[95:80])
  );


  bsg_mux_one_hot_width_p16_els_p16
  \l_6_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[111:96]),
    .data_o(o[111:96])
  );


  bsg_mux_one_hot_width_p16_els_p16
  \l_7_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[127:112]),
    .data_o(o[127:112])
  );


  bsg_mux_one_hot_width_p16_els_p16
  \l_8_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[143:128]),
    .data_o(o[143:128])
  );


  bsg_mux_one_hot_width_p16_els_p16
  \l_9_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[159:144]),
    .data_o(o[159:144])
  );


  bsg_mux_one_hot_width_p16_els_p16
  \l_10_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[175:160]),
    .data_o(o[175:160])
  );


  bsg_mux_one_hot_width_p16_els_p16
  \l_11_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[191:176]),
    .data_o(o[191:176])
  );


  bsg_mux_one_hot_width_p16_els_p16
  \l_12_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[207:192]),
    .data_o(o[207:192])
  );


  bsg_mux_one_hot_width_p16_els_p16
  \l_13_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[223:208]),
    .data_o(o[223:208])
  );


  bsg_mux_one_hot_width_p16_els_p16
  \l_14_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[239:224]),
    .data_o(o[239:224])
  );


  bsg_mux_one_hot_width_p16_els_p16
  \l_15_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[255:240]),
    .data_o(o[255:240])
  );


endmodule

