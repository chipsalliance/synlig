

module top
(
  clk_i,
  reset_i,
  valid_i,
  data_i,
  ready_o,
  valid_o,
  data_o,
  yumi_cnt_i
);

  input [15:0] data_i;
  output [31:0] valid_o;
  output [511:0] data_o;
  input [5:0] yumi_cnt_i;
  input clk_i;
  input reset_i;
  input valid_i;
  output ready_o;

  bsg_serial_in_parallel_out
  wrapper
  (
    .data_i(data_i),
    .valid_o(valid_o),
    .data_o(data_o),
    .yumi_cnt_i(yumi_cnt_i),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .valid_i(valid_i),
    .ready_o(ready_o)
  );


endmodule



module bsg_serial_in_parallel_out
(
  clk_i,
  reset_i,
  valid_i,
  data_i,
  ready_o,
  valid_o,
  data_o,
  yumi_cnt_i
);

  input [15:0] data_i;
  output [31:0] valid_o;
  output [511:0] data_o;
  input [5:0] yumi_cnt_i;
  input clk_i;
  input reset_i;
  input valid_i;
  output ready_o;
  wire [31:0] valid_o,valid_r,valid_nn;
  wire [511:0] data_o,data_r,data_nn;
  wire ready_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
  N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,
  N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,
  N404,N405,N406,N407,N408,data_n_63__15_,data_n_63__14_,data_n_63__13_,
  data_n_63__12_,data_n_63__11_,data_n_63__10_,data_n_63__9_,data_n_63__8_,data_n_63__7_,
  data_n_63__6_,data_n_63__5_,data_n_63__4_,data_n_63__3_,data_n_63__2_,data_n_63__1_,
  data_n_63__0_,data_n_62__15_,data_n_62__14_,data_n_62__13_,data_n_62__12_,
  data_n_62__11_,data_n_62__10_,data_n_62__9_,data_n_62__8_,data_n_62__7_,data_n_62__6_,
  data_n_62__5_,data_n_62__4_,data_n_62__3_,data_n_62__2_,data_n_62__1_,
  data_n_62__0_,data_n_61__15_,data_n_61__14_,data_n_61__13_,data_n_61__12_,data_n_61__11_,
  data_n_61__10_,data_n_61__9_,data_n_61__8_,data_n_61__7_,data_n_61__6_,
  data_n_61__5_,data_n_61__4_,data_n_61__3_,data_n_61__2_,data_n_61__1_,data_n_61__0_,
  data_n_60__15_,data_n_60__14_,data_n_60__13_,data_n_60__12_,data_n_60__11_,
  data_n_60__10_,data_n_60__9_,data_n_60__8_,data_n_60__7_,data_n_60__6_,data_n_60__5_,
  data_n_60__4_,data_n_60__3_,data_n_60__2_,data_n_60__1_,data_n_60__0_,data_n_59__15_,
  data_n_59__14_,data_n_59__13_,data_n_59__12_,data_n_59__11_,data_n_59__10_,
  data_n_59__9_,data_n_59__8_,data_n_59__7_,data_n_59__6_,data_n_59__5_,data_n_59__4_,
  data_n_59__3_,data_n_59__2_,data_n_59__1_,data_n_59__0_,data_n_58__15_,
  data_n_58__14_,data_n_58__13_,data_n_58__12_,data_n_58__11_,data_n_58__10_,data_n_58__9_,
  data_n_58__8_,data_n_58__7_,data_n_58__6_,data_n_58__5_,data_n_58__4_,
  data_n_58__3_,data_n_58__2_,data_n_58__1_,data_n_58__0_,data_n_57__15_,data_n_57__14_,
  data_n_57__13_,data_n_57__12_,data_n_57__11_,data_n_57__10_,data_n_57__9_,
  data_n_57__8_,data_n_57__7_,data_n_57__6_,data_n_57__5_,data_n_57__4_,data_n_57__3_,
  data_n_57__2_,data_n_57__1_,data_n_57__0_,data_n_56__15_,data_n_56__14_,data_n_56__13_,
  data_n_56__12_,data_n_56__11_,data_n_56__10_,data_n_56__9_,data_n_56__8_,
  data_n_56__7_,data_n_56__6_,data_n_56__5_,data_n_56__4_,data_n_56__3_,data_n_56__2_,
  data_n_56__1_,data_n_56__0_,data_n_55__15_,data_n_55__14_,data_n_55__13_,
  data_n_55__12_,data_n_55__11_,data_n_55__10_,data_n_55__9_,data_n_55__8_,data_n_55__7_,
  data_n_55__6_,data_n_55__5_,data_n_55__4_,data_n_55__3_,data_n_55__2_,data_n_55__1_,
  data_n_55__0_,data_n_54__15_,data_n_54__14_,data_n_54__13_,data_n_54__12_,
  data_n_54__11_,data_n_54__10_,data_n_54__9_,data_n_54__8_,data_n_54__7_,data_n_54__6_,
  data_n_54__5_,data_n_54__4_,data_n_54__3_,data_n_54__2_,data_n_54__1_,
  data_n_54__0_,data_n_53__15_,data_n_53__14_,data_n_53__13_,data_n_53__12_,data_n_53__11_,
  data_n_53__10_,data_n_53__9_,data_n_53__8_,data_n_53__7_,data_n_53__6_,
  data_n_53__5_,data_n_53__4_,data_n_53__3_,data_n_53__2_,data_n_53__1_,data_n_53__0_,
  data_n_52__15_,data_n_52__14_,data_n_52__13_,data_n_52__12_,data_n_52__11_,
  data_n_52__10_,data_n_52__9_,data_n_52__8_,data_n_52__7_,data_n_52__6_,data_n_52__5_,
  data_n_52__4_,data_n_52__3_,data_n_52__2_,data_n_52__1_,data_n_52__0_,data_n_51__15_,
  data_n_51__14_,data_n_51__13_,data_n_51__12_,data_n_51__11_,data_n_51__10_,
  data_n_51__9_,data_n_51__8_,data_n_51__7_,data_n_51__6_,data_n_51__5_,data_n_51__4_,
  data_n_51__3_,data_n_51__2_,data_n_51__1_,data_n_51__0_,data_n_50__15_,
  data_n_50__14_,data_n_50__13_,data_n_50__12_,data_n_50__11_,data_n_50__10_,data_n_50__9_,
  data_n_50__8_,data_n_50__7_,data_n_50__6_,data_n_50__5_,data_n_50__4_,
  data_n_50__3_,data_n_50__2_,data_n_50__1_,data_n_50__0_,data_n_49__15_,data_n_49__14_,
  data_n_49__13_,data_n_49__12_,data_n_49__11_,data_n_49__10_,data_n_49__9_,
  data_n_49__8_,data_n_49__7_,data_n_49__6_,data_n_49__5_,data_n_49__4_,data_n_49__3_,
  data_n_49__2_,data_n_49__1_,data_n_49__0_,data_n_48__15_,data_n_48__14_,data_n_48__13_,
  data_n_48__12_,data_n_48__11_,data_n_48__10_,data_n_48__9_,data_n_48__8_,
  data_n_48__7_,data_n_48__6_,data_n_48__5_,data_n_48__4_,data_n_48__3_,data_n_48__2_,
  data_n_48__1_,data_n_48__0_,data_n_47__15_,data_n_47__14_,data_n_47__13_,
  data_n_47__12_,data_n_47__11_,data_n_47__10_,data_n_47__9_,data_n_47__8_,data_n_47__7_,
  data_n_47__6_,data_n_47__5_,data_n_47__4_,data_n_47__3_,data_n_47__2_,data_n_47__1_,
  data_n_47__0_,data_n_46__15_,data_n_46__14_,data_n_46__13_,data_n_46__12_,
  data_n_46__11_,data_n_46__10_,data_n_46__9_,data_n_46__8_,data_n_46__7_,data_n_46__6_,
  data_n_46__5_,data_n_46__4_,data_n_46__3_,data_n_46__2_,data_n_46__1_,
  data_n_46__0_,data_n_45__15_,data_n_45__14_,data_n_45__13_,data_n_45__12_,data_n_45__11_,
  data_n_45__10_,data_n_45__9_,data_n_45__8_,data_n_45__7_,data_n_45__6_,
  data_n_45__5_,data_n_45__4_,data_n_45__3_,data_n_45__2_,data_n_45__1_,data_n_45__0_,
  data_n_44__15_,data_n_44__14_,data_n_44__13_,data_n_44__12_,data_n_44__11_,
  data_n_44__10_,data_n_44__9_,data_n_44__8_,data_n_44__7_,data_n_44__6_,data_n_44__5_,
  data_n_44__4_,data_n_44__3_,data_n_44__2_,data_n_44__1_,data_n_44__0_,data_n_43__15_,
  data_n_43__14_,data_n_43__13_,data_n_43__12_,data_n_43__11_,data_n_43__10_,
  data_n_43__9_,data_n_43__8_,data_n_43__7_,data_n_43__6_,data_n_43__5_,data_n_43__4_,
  data_n_43__3_,data_n_43__2_,data_n_43__1_,data_n_43__0_,data_n_42__15_,
  data_n_42__14_,data_n_42__13_,data_n_42__12_,data_n_42__11_,data_n_42__10_,data_n_42__9_,
  data_n_42__8_,data_n_42__7_,data_n_42__6_,data_n_42__5_,data_n_42__4_,
  data_n_42__3_,data_n_42__2_,data_n_42__1_,data_n_42__0_,data_n_41__15_,data_n_41__14_,
  data_n_41__13_,data_n_41__12_,data_n_41__11_,data_n_41__10_,data_n_41__9_,
  data_n_41__8_,data_n_41__7_,data_n_41__6_,data_n_41__5_,data_n_41__4_,data_n_41__3_,
  data_n_41__2_,data_n_41__1_,data_n_41__0_,data_n_40__15_,data_n_40__14_,data_n_40__13_,
  data_n_40__12_,data_n_40__11_,data_n_40__10_,data_n_40__9_,data_n_40__8_,
  data_n_40__7_,data_n_40__6_,data_n_40__5_,data_n_40__4_,data_n_40__3_,data_n_40__2_,
  data_n_40__1_,data_n_40__0_,data_n_39__15_,data_n_39__14_,data_n_39__13_,
  data_n_39__12_,data_n_39__11_,data_n_39__10_,data_n_39__9_,data_n_39__8_,data_n_39__7_,
  data_n_39__6_,data_n_39__5_,data_n_39__4_,data_n_39__3_,data_n_39__2_,data_n_39__1_,
  data_n_39__0_,data_n_38__15_,data_n_38__14_,data_n_38__13_,data_n_38__12_,
  data_n_38__11_,data_n_38__10_,data_n_38__9_,data_n_38__8_,data_n_38__7_,data_n_38__6_,
  data_n_38__5_,data_n_38__4_,data_n_38__3_,data_n_38__2_,data_n_38__1_,
  data_n_38__0_,data_n_37__15_,data_n_37__14_,data_n_37__13_,data_n_37__12_,data_n_37__11_,
  data_n_37__10_,data_n_37__9_,data_n_37__8_,data_n_37__7_,data_n_37__6_,
  data_n_37__5_,data_n_37__4_,data_n_37__3_,data_n_37__2_,data_n_37__1_,data_n_37__0_,
  data_n_36__15_,data_n_36__14_,data_n_36__13_,data_n_36__12_,data_n_36__11_,
  data_n_36__10_,data_n_36__9_,data_n_36__8_,data_n_36__7_,data_n_36__6_,data_n_36__5_,
  data_n_36__4_,data_n_36__3_,data_n_36__2_,data_n_36__1_,data_n_36__0_,data_n_35__15_,
  data_n_35__14_,data_n_35__13_,data_n_35__12_,data_n_35__11_,data_n_35__10_,
  data_n_35__9_,data_n_35__8_,data_n_35__7_,data_n_35__6_,data_n_35__5_,data_n_35__4_,
  data_n_35__3_,data_n_35__2_,data_n_35__1_,data_n_35__0_,data_n_34__15_,
  data_n_34__14_,data_n_34__13_,data_n_34__12_,data_n_34__11_,data_n_34__10_,data_n_34__9_,
  data_n_34__8_,data_n_34__7_,data_n_34__6_,data_n_34__5_,data_n_34__4_,
  data_n_34__3_,data_n_34__2_,data_n_34__1_,data_n_34__0_,data_n_33__15_,data_n_33__14_,
  data_n_33__13_,data_n_33__12_,data_n_33__11_,data_n_33__10_,data_n_33__9_,
  data_n_33__8_,data_n_33__7_,data_n_33__6_,data_n_33__5_,data_n_33__4_,data_n_33__3_,
  data_n_33__2_,data_n_33__1_,data_n_33__0_,data_n_32__15_,data_n_32__14_,data_n_32__13_,
  data_n_32__12_,data_n_32__11_,data_n_32__10_,data_n_32__9_,data_n_32__8_,
  data_n_32__7_,data_n_32__6_,data_n_32__5_,data_n_32__4_,data_n_32__3_,data_n_32__2_,
  data_n_32__1_,data_n_32__0_,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,
  N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,
  N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,
  N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,
  N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,
  N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,
  N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,
  N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,
  N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,
  N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
  N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,
  N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,
  N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,
  N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,
  N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,
  N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,
  N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,
  N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,
  N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,
  N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,
  N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,
  N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,
  N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,
  N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,
  N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,
  N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,
  N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,
  N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,
  N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,
  N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,
  N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
  N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,
  N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,
  N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,
  N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,
  N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,
  N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,
  N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,
  N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,
  N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,
  N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,
  N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,
  N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,
  N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,
  N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,
  N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,
  N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,
  N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,
  N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,
  N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,
  N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,
  N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,
  N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,
  N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,
  N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,
  N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,
  N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,
  N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,
  N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,
  N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,
  N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
  N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,
  N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,
  N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,
  N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369;
  wire [5:0] num_els_r,num_els_n;
  wire [63:32] valid_n;
  reg valid_r_31_sv2v_reg,valid_r_30_sv2v_reg,valid_r_29_sv2v_reg,valid_r_28_sv2v_reg,
  valid_r_27_sv2v_reg,valid_r_26_sv2v_reg,valid_r_25_sv2v_reg,valid_r_24_sv2v_reg,
  valid_r_23_sv2v_reg,valid_r_22_sv2v_reg,valid_r_21_sv2v_reg,valid_r_20_sv2v_reg,
  valid_r_19_sv2v_reg,valid_r_18_sv2v_reg,valid_r_17_sv2v_reg,valid_r_16_sv2v_reg,
  valid_r_15_sv2v_reg,valid_r_14_sv2v_reg,valid_r_13_sv2v_reg,valid_r_12_sv2v_reg,
  valid_r_11_sv2v_reg,valid_r_10_sv2v_reg,valid_r_9_sv2v_reg,valid_r_8_sv2v_reg,
  valid_r_7_sv2v_reg,valid_r_6_sv2v_reg,valid_r_5_sv2v_reg,valid_r_4_sv2v_reg,
  valid_r_3_sv2v_reg,valid_r_2_sv2v_reg,valid_r_1_sv2v_reg,valid_r_0_sv2v_reg,
  num_els_r_5_sv2v_reg,num_els_r_4_sv2v_reg,num_els_r_3_sv2v_reg,num_els_r_2_sv2v_reg,
  num_els_r_1_sv2v_reg,num_els_r_0_sv2v_reg,data_r_511_sv2v_reg,data_r_510_sv2v_reg,
  data_r_509_sv2v_reg,data_r_508_sv2v_reg,data_r_507_sv2v_reg,data_r_506_sv2v_reg,
  data_r_505_sv2v_reg,data_r_504_sv2v_reg,data_r_503_sv2v_reg,data_r_502_sv2v_reg,
  data_r_501_sv2v_reg,data_r_500_sv2v_reg,data_r_499_sv2v_reg,data_r_498_sv2v_reg,
  data_r_497_sv2v_reg,data_r_496_sv2v_reg,data_r_495_sv2v_reg,data_r_494_sv2v_reg,
  data_r_493_sv2v_reg,data_r_492_sv2v_reg,data_r_491_sv2v_reg,data_r_490_sv2v_reg,
  data_r_489_sv2v_reg,data_r_488_sv2v_reg,data_r_487_sv2v_reg,data_r_486_sv2v_reg,
  data_r_485_sv2v_reg,data_r_484_sv2v_reg,data_r_483_sv2v_reg,data_r_482_sv2v_reg,
  data_r_481_sv2v_reg,data_r_480_sv2v_reg,data_r_479_sv2v_reg,data_r_478_sv2v_reg,
  data_r_477_sv2v_reg,data_r_476_sv2v_reg,data_r_475_sv2v_reg,data_r_474_sv2v_reg,
  data_r_473_sv2v_reg,data_r_472_sv2v_reg,data_r_471_sv2v_reg,data_r_470_sv2v_reg,
  data_r_469_sv2v_reg,data_r_468_sv2v_reg,data_r_467_sv2v_reg,data_r_466_sv2v_reg,
  data_r_465_sv2v_reg,data_r_464_sv2v_reg,data_r_463_sv2v_reg,data_r_462_sv2v_reg,
  data_r_461_sv2v_reg,data_r_460_sv2v_reg,data_r_459_sv2v_reg,data_r_458_sv2v_reg,
  data_r_457_sv2v_reg,data_r_456_sv2v_reg,data_r_455_sv2v_reg,data_r_454_sv2v_reg,
  data_r_453_sv2v_reg,data_r_452_sv2v_reg,data_r_451_sv2v_reg,data_r_450_sv2v_reg,
  data_r_449_sv2v_reg,data_r_448_sv2v_reg,data_r_447_sv2v_reg,data_r_446_sv2v_reg,
  data_r_445_sv2v_reg,data_r_444_sv2v_reg,data_r_443_sv2v_reg,data_r_442_sv2v_reg,
  data_r_441_sv2v_reg,data_r_440_sv2v_reg,data_r_439_sv2v_reg,data_r_438_sv2v_reg,
  data_r_437_sv2v_reg,data_r_436_sv2v_reg,data_r_435_sv2v_reg,data_r_434_sv2v_reg,
  data_r_433_sv2v_reg,data_r_432_sv2v_reg,data_r_431_sv2v_reg,data_r_430_sv2v_reg,
  data_r_429_sv2v_reg,data_r_428_sv2v_reg,data_r_427_sv2v_reg,data_r_426_sv2v_reg,
  data_r_425_sv2v_reg,data_r_424_sv2v_reg,data_r_423_sv2v_reg,data_r_422_sv2v_reg,
  data_r_421_sv2v_reg,data_r_420_sv2v_reg,data_r_419_sv2v_reg,data_r_418_sv2v_reg,
  data_r_417_sv2v_reg,data_r_416_sv2v_reg,data_r_415_sv2v_reg,data_r_414_sv2v_reg,
  data_r_413_sv2v_reg,data_r_412_sv2v_reg,data_r_411_sv2v_reg,data_r_410_sv2v_reg,
  data_r_409_sv2v_reg,data_r_408_sv2v_reg,data_r_407_sv2v_reg,data_r_406_sv2v_reg,
  data_r_405_sv2v_reg,data_r_404_sv2v_reg,data_r_403_sv2v_reg,data_r_402_sv2v_reg,
  data_r_401_sv2v_reg,data_r_400_sv2v_reg,data_r_399_sv2v_reg,data_r_398_sv2v_reg,
  data_r_397_sv2v_reg,data_r_396_sv2v_reg,data_r_395_sv2v_reg,data_r_394_sv2v_reg,
  data_r_393_sv2v_reg,data_r_392_sv2v_reg,data_r_391_sv2v_reg,data_r_390_sv2v_reg,
  data_r_389_sv2v_reg,data_r_388_sv2v_reg,data_r_387_sv2v_reg,data_r_386_sv2v_reg,
  data_r_385_sv2v_reg,data_r_384_sv2v_reg,data_r_383_sv2v_reg,data_r_382_sv2v_reg,
  data_r_381_sv2v_reg,data_r_380_sv2v_reg,data_r_379_sv2v_reg,data_r_378_sv2v_reg,
  data_r_377_sv2v_reg,data_r_376_sv2v_reg,data_r_375_sv2v_reg,data_r_374_sv2v_reg,
  data_r_373_sv2v_reg,data_r_372_sv2v_reg,data_r_371_sv2v_reg,data_r_370_sv2v_reg,
  data_r_369_sv2v_reg,data_r_368_sv2v_reg,data_r_367_sv2v_reg,data_r_366_sv2v_reg,
  data_r_365_sv2v_reg,data_r_364_sv2v_reg,data_r_363_sv2v_reg,data_r_362_sv2v_reg,
  data_r_361_sv2v_reg,data_r_360_sv2v_reg,data_r_359_sv2v_reg,data_r_358_sv2v_reg,
  data_r_357_sv2v_reg,data_r_356_sv2v_reg,data_r_355_sv2v_reg,data_r_354_sv2v_reg,
  data_r_353_sv2v_reg,data_r_352_sv2v_reg,data_r_351_sv2v_reg,data_r_350_sv2v_reg,
  data_r_349_sv2v_reg,data_r_348_sv2v_reg,data_r_347_sv2v_reg,data_r_346_sv2v_reg,
  data_r_345_sv2v_reg,data_r_344_sv2v_reg,data_r_343_sv2v_reg,data_r_342_sv2v_reg,
  data_r_341_sv2v_reg,data_r_340_sv2v_reg,data_r_339_sv2v_reg,data_r_338_sv2v_reg,
  data_r_337_sv2v_reg,data_r_336_sv2v_reg,data_r_335_sv2v_reg,data_r_334_sv2v_reg,
  data_r_333_sv2v_reg,data_r_332_sv2v_reg,data_r_331_sv2v_reg,data_r_330_sv2v_reg,
  data_r_329_sv2v_reg,data_r_328_sv2v_reg,data_r_327_sv2v_reg,data_r_326_sv2v_reg,
  data_r_325_sv2v_reg,data_r_324_sv2v_reg,data_r_323_sv2v_reg,data_r_322_sv2v_reg,
  data_r_321_sv2v_reg,data_r_320_sv2v_reg,data_r_319_sv2v_reg,data_r_318_sv2v_reg,
  data_r_317_sv2v_reg,data_r_316_sv2v_reg,data_r_315_sv2v_reg,data_r_314_sv2v_reg,
  data_r_313_sv2v_reg,data_r_312_sv2v_reg,data_r_311_sv2v_reg,data_r_310_sv2v_reg,
  data_r_309_sv2v_reg,data_r_308_sv2v_reg,data_r_307_sv2v_reg,data_r_306_sv2v_reg,
  data_r_305_sv2v_reg,data_r_304_sv2v_reg,data_r_303_sv2v_reg,data_r_302_sv2v_reg,
  data_r_301_sv2v_reg,data_r_300_sv2v_reg,data_r_299_sv2v_reg,data_r_298_sv2v_reg,
  data_r_297_sv2v_reg,data_r_296_sv2v_reg,data_r_295_sv2v_reg,data_r_294_sv2v_reg,
  data_r_293_sv2v_reg,data_r_292_sv2v_reg,data_r_291_sv2v_reg,data_r_290_sv2v_reg,
  data_r_289_sv2v_reg,data_r_288_sv2v_reg,data_r_287_sv2v_reg,data_r_286_sv2v_reg,
  data_r_285_sv2v_reg,data_r_284_sv2v_reg,data_r_283_sv2v_reg,data_r_282_sv2v_reg,
  data_r_281_sv2v_reg,data_r_280_sv2v_reg,data_r_279_sv2v_reg,data_r_278_sv2v_reg,
  data_r_277_sv2v_reg,data_r_276_sv2v_reg,data_r_275_sv2v_reg,data_r_274_sv2v_reg,
  data_r_273_sv2v_reg,data_r_272_sv2v_reg,data_r_271_sv2v_reg,data_r_270_sv2v_reg,
  data_r_269_sv2v_reg,data_r_268_sv2v_reg,data_r_267_sv2v_reg,data_r_266_sv2v_reg,
  data_r_265_sv2v_reg,data_r_264_sv2v_reg,data_r_263_sv2v_reg,data_r_262_sv2v_reg,
  data_r_261_sv2v_reg,data_r_260_sv2v_reg,data_r_259_sv2v_reg,data_r_258_sv2v_reg,
  data_r_257_sv2v_reg,data_r_256_sv2v_reg,data_r_255_sv2v_reg,data_r_254_sv2v_reg,
  data_r_253_sv2v_reg,data_r_252_sv2v_reg,data_r_251_sv2v_reg,data_r_250_sv2v_reg,
  data_r_249_sv2v_reg,data_r_248_sv2v_reg,data_r_247_sv2v_reg,data_r_246_sv2v_reg,
  data_r_245_sv2v_reg,data_r_244_sv2v_reg,data_r_243_sv2v_reg,data_r_242_sv2v_reg,
  data_r_241_sv2v_reg,data_r_240_sv2v_reg,data_r_239_sv2v_reg,data_r_238_sv2v_reg,
  data_r_237_sv2v_reg,data_r_236_sv2v_reg,data_r_235_sv2v_reg,data_r_234_sv2v_reg,
  data_r_233_sv2v_reg,data_r_232_sv2v_reg,data_r_231_sv2v_reg,data_r_230_sv2v_reg,
  data_r_229_sv2v_reg,data_r_228_sv2v_reg,data_r_227_sv2v_reg,data_r_226_sv2v_reg,
  data_r_225_sv2v_reg,data_r_224_sv2v_reg,data_r_223_sv2v_reg,data_r_222_sv2v_reg,
  data_r_221_sv2v_reg,data_r_220_sv2v_reg,data_r_219_sv2v_reg,data_r_218_sv2v_reg,
  data_r_217_sv2v_reg,data_r_216_sv2v_reg,data_r_215_sv2v_reg,data_r_214_sv2v_reg,
  data_r_213_sv2v_reg,data_r_212_sv2v_reg,data_r_211_sv2v_reg,data_r_210_sv2v_reg,
  data_r_209_sv2v_reg,data_r_208_sv2v_reg,data_r_207_sv2v_reg,data_r_206_sv2v_reg,
  data_r_205_sv2v_reg,data_r_204_sv2v_reg,data_r_203_sv2v_reg,data_r_202_sv2v_reg,
  data_r_201_sv2v_reg,data_r_200_sv2v_reg,data_r_199_sv2v_reg,data_r_198_sv2v_reg,
  data_r_197_sv2v_reg,data_r_196_sv2v_reg,data_r_195_sv2v_reg,data_r_194_sv2v_reg,
  data_r_193_sv2v_reg,data_r_192_sv2v_reg,data_r_191_sv2v_reg,data_r_190_sv2v_reg,
  data_r_189_sv2v_reg,data_r_188_sv2v_reg,data_r_187_sv2v_reg,data_r_186_sv2v_reg,
  data_r_185_sv2v_reg,data_r_184_sv2v_reg,data_r_183_sv2v_reg,data_r_182_sv2v_reg,
  data_r_181_sv2v_reg,data_r_180_sv2v_reg,data_r_179_sv2v_reg,data_r_178_sv2v_reg,
  data_r_177_sv2v_reg,data_r_176_sv2v_reg,data_r_175_sv2v_reg,data_r_174_sv2v_reg,
  data_r_173_sv2v_reg,data_r_172_sv2v_reg,data_r_171_sv2v_reg,data_r_170_sv2v_reg,
  data_r_169_sv2v_reg,data_r_168_sv2v_reg,data_r_167_sv2v_reg,data_r_166_sv2v_reg,
  data_r_165_sv2v_reg,data_r_164_sv2v_reg,data_r_163_sv2v_reg,data_r_162_sv2v_reg,
  data_r_161_sv2v_reg,data_r_160_sv2v_reg,data_r_159_sv2v_reg,data_r_158_sv2v_reg,
  data_r_157_sv2v_reg,data_r_156_sv2v_reg,data_r_155_sv2v_reg,data_r_154_sv2v_reg,
  data_r_153_sv2v_reg,data_r_152_sv2v_reg,data_r_151_sv2v_reg,data_r_150_sv2v_reg,
  data_r_149_sv2v_reg,data_r_148_sv2v_reg,data_r_147_sv2v_reg,data_r_146_sv2v_reg,
  data_r_145_sv2v_reg,data_r_144_sv2v_reg,data_r_143_sv2v_reg,data_r_142_sv2v_reg,
  data_r_141_sv2v_reg,data_r_140_sv2v_reg,data_r_139_sv2v_reg,data_r_138_sv2v_reg,
  data_r_137_sv2v_reg,data_r_136_sv2v_reg,data_r_135_sv2v_reg,data_r_134_sv2v_reg,
  data_r_133_sv2v_reg,data_r_132_sv2v_reg,data_r_131_sv2v_reg,data_r_130_sv2v_reg,
  data_r_129_sv2v_reg,data_r_128_sv2v_reg,data_r_127_sv2v_reg,data_r_126_sv2v_reg,
  data_r_125_sv2v_reg,data_r_124_sv2v_reg,data_r_123_sv2v_reg,data_r_122_sv2v_reg,
  data_r_121_sv2v_reg,data_r_120_sv2v_reg,data_r_119_sv2v_reg,data_r_118_sv2v_reg,
  data_r_117_sv2v_reg,data_r_116_sv2v_reg,data_r_115_sv2v_reg,data_r_114_sv2v_reg,
  data_r_113_sv2v_reg,data_r_112_sv2v_reg,data_r_111_sv2v_reg,data_r_110_sv2v_reg,
  data_r_109_sv2v_reg,data_r_108_sv2v_reg,data_r_107_sv2v_reg,data_r_106_sv2v_reg,
  data_r_105_sv2v_reg,data_r_104_sv2v_reg,data_r_103_sv2v_reg,data_r_102_sv2v_reg,
  data_r_101_sv2v_reg,data_r_100_sv2v_reg,data_r_99_sv2v_reg,data_r_98_sv2v_reg,
  data_r_97_sv2v_reg,data_r_96_sv2v_reg,data_r_95_sv2v_reg,data_r_94_sv2v_reg,
  data_r_93_sv2v_reg,data_r_92_sv2v_reg,data_r_91_sv2v_reg,data_r_90_sv2v_reg,
  data_r_89_sv2v_reg,data_r_88_sv2v_reg,data_r_87_sv2v_reg,data_r_86_sv2v_reg,
  data_r_85_sv2v_reg,data_r_84_sv2v_reg,data_r_83_sv2v_reg,data_r_82_sv2v_reg,data_r_81_sv2v_reg,
  data_r_80_sv2v_reg,data_r_79_sv2v_reg,data_r_78_sv2v_reg,data_r_77_sv2v_reg,
  data_r_76_sv2v_reg,data_r_75_sv2v_reg,data_r_74_sv2v_reg,data_r_73_sv2v_reg,
  data_r_72_sv2v_reg,data_r_71_sv2v_reg,data_r_70_sv2v_reg,data_r_69_sv2v_reg,
  data_r_68_sv2v_reg,data_r_67_sv2v_reg,data_r_66_sv2v_reg,data_r_65_sv2v_reg,data_r_64_sv2v_reg,
  data_r_63_sv2v_reg,data_r_62_sv2v_reg,data_r_61_sv2v_reg,data_r_60_sv2v_reg,
  data_r_59_sv2v_reg,data_r_58_sv2v_reg,data_r_57_sv2v_reg,data_r_56_sv2v_reg,
  data_r_55_sv2v_reg,data_r_54_sv2v_reg,data_r_53_sv2v_reg,data_r_52_sv2v_reg,
  data_r_51_sv2v_reg,data_r_50_sv2v_reg,data_r_49_sv2v_reg,data_r_48_sv2v_reg,
  data_r_47_sv2v_reg,data_r_46_sv2v_reg,data_r_45_sv2v_reg,data_r_44_sv2v_reg,data_r_43_sv2v_reg,
  data_r_42_sv2v_reg,data_r_41_sv2v_reg,data_r_40_sv2v_reg,data_r_39_sv2v_reg,
  data_r_38_sv2v_reg,data_r_37_sv2v_reg,data_r_36_sv2v_reg,data_r_35_sv2v_reg,
  data_r_34_sv2v_reg,data_r_33_sv2v_reg,data_r_32_sv2v_reg,data_r_31_sv2v_reg,
  data_r_30_sv2v_reg,data_r_29_sv2v_reg,data_r_28_sv2v_reg,data_r_27_sv2v_reg,
  data_r_26_sv2v_reg,data_r_25_sv2v_reg,data_r_24_sv2v_reg,data_r_23_sv2v_reg,data_r_22_sv2v_reg,
  data_r_21_sv2v_reg,data_r_20_sv2v_reg,data_r_19_sv2v_reg,data_r_18_sv2v_reg,
  data_r_17_sv2v_reg,data_r_16_sv2v_reg,data_r_15_sv2v_reg,data_r_14_sv2v_reg,
  data_r_13_sv2v_reg,data_r_12_sv2v_reg,data_r_11_sv2v_reg,data_r_10_sv2v_reg,
  data_r_9_sv2v_reg,data_r_8_sv2v_reg,data_r_7_sv2v_reg,data_r_6_sv2v_reg,data_r_5_sv2v_reg,
  data_r_4_sv2v_reg,data_r_3_sv2v_reg,data_r_2_sv2v_reg,data_r_1_sv2v_reg,
  data_r_0_sv2v_reg;
  assign valid_r[31] = valid_r_31_sv2v_reg;
  assign valid_r[30] = valid_r_30_sv2v_reg;
  assign valid_r[29] = valid_r_29_sv2v_reg;
  assign valid_r[28] = valid_r_28_sv2v_reg;
  assign valid_r[27] = valid_r_27_sv2v_reg;
  assign valid_r[26] = valid_r_26_sv2v_reg;
  assign valid_r[25] = valid_r_25_sv2v_reg;
  assign valid_r[24] = valid_r_24_sv2v_reg;
  assign valid_r[23] = valid_r_23_sv2v_reg;
  assign valid_r[22] = valid_r_22_sv2v_reg;
  assign valid_r[21] = valid_r_21_sv2v_reg;
  assign valid_r[20] = valid_r_20_sv2v_reg;
  assign valid_r[19] = valid_r_19_sv2v_reg;
  assign valid_r[18] = valid_r_18_sv2v_reg;
  assign valid_r[17] = valid_r_17_sv2v_reg;
  assign valid_r[16] = valid_r_16_sv2v_reg;
  assign valid_r[15] = valid_r_15_sv2v_reg;
  assign valid_r[14] = valid_r_14_sv2v_reg;
  assign valid_r[13] = valid_r_13_sv2v_reg;
  assign valid_r[12] = valid_r_12_sv2v_reg;
  assign valid_r[11] = valid_r_11_sv2v_reg;
  assign valid_r[10] = valid_r_10_sv2v_reg;
  assign valid_r[9] = valid_r_9_sv2v_reg;
  assign valid_r[8] = valid_r_8_sv2v_reg;
  assign valid_r[7] = valid_r_7_sv2v_reg;
  assign valid_r[6] = valid_r_6_sv2v_reg;
  assign valid_r[5] = valid_r_5_sv2v_reg;
  assign valid_r[4] = valid_r_4_sv2v_reg;
  assign valid_r[3] = valid_r_3_sv2v_reg;
  assign valid_r[2] = valid_r_2_sv2v_reg;
  assign valid_r[1] = valid_r_1_sv2v_reg;
  assign valid_r[0] = valid_r_0_sv2v_reg;
  assign num_els_r[5] = num_els_r_5_sv2v_reg;
  assign num_els_r[4] = num_els_r_4_sv2v_reg;
  assign num_els_r[3] = num_els_r_3_sv2v_reg;
  assign num_els_r[2] = num_els_r_2_sv2v_reg;
  assign num_els_r[1] = num_els_r_1_sv2v_reg;
  assign num_els_r[0] = num_els_r_0_sv2v_reg;
  assign data_r[511] = data_r_511_sv2v_reg;
  assign data_r[510] = data_r_510_sv2v_reg;
  assign data_r[509] = data_r_509_sv2v_reg;
  assign data_r[508] = data_r_508_sv2v_reg;
  assign data_r[507] = data_r_507_sv2v_reg;
  assign data_r[506] = data_r_506_sv2v_reg;
  assign data_r[505] = data_r_505_sv2v_reg;
  assign data_r[504] = data_r_504_sv2v_reg;
  assign data_r[503] = data_r_503_sv2v_reg;
  assign data_r[502] = data_r_502_sv2v_reg;
  assign data_r[501] = data_r_501_sv2v_reg;
  assign data_r[500] = data_r_500_sv2v_reg;
  assign data_r[499] = data_r_499_sv2v_reg;
  assign data_r[498] = data_r_498_sv2v_reg;
  assign data_r[497] = data_r_497_sv2v_reg;
  assign data_r[496] = data_r_496_sv2v_reg;
  assign data_r[495] = data_r_495_sv2v_reg;
  assign data_r[494] = data_r_494_sv2v_reg;
  assign data_r[493] = data_r_493_sv2v_reg;
  assign data_r[492] = data_r_492_sv2v_reg;
  assign data_r[491] = data_r_491_sv2v_reg;
  assign data_r[490] = data_r_490_sv2v_reg;
  assign data_r[489] = data_r_489_sv2v_reg;
  assign data_r[488] = data_r_488_sv2v_reg;
  assign data_r[487] = data_r_487_sv2v_reg;
  assign data_r[486] = data_r_486_sv2v_reg;
  assign data_r[485] = data_r_485_sv2v_reg;
  assign data_r[484] = data_r_484_sv2v_reg;
  assign data_r[483] = data_r_483_sv2v_reg;
  assign data_r[482] = data_r_482_sv2v_reg;
  assign data_r[481] = data_r_481_sv2v_reg;
  assign data_r[480] = data_r_480_sv2v_reg;
  assign data_r[479] = data_r_479_sv2v_reg;
  assign data_r[478] = data_r_478_sv2v_reg;
  assign data_r[477] = data_r_477_sv2v_reg;
  assign data_r[476] = data_r_476_sv2v_reg;
  assign data_r[475] = data_r_475_sv2v_reg;
  assign data_r[474] = data_r_474_sv2v_reg;
  assign data_r[473] = data_r_473_sv2v_reg;
  assign data_r[472] = data_r_472_sv2v_reg;
  assign data_r[471] = data_r_471_sv2v_reg;
  assign data_r[470] = data_r_470_sv2v_reg;
  assign data_r[469] = data_r_469_sv2v_reg;
  assign data_r[468] = data_r_468_sv2v_reg;
  assign data_r[467] = data_r_467_sv2v_reg;
  assign data_r[466] = data_r_466_sv2v_reg;
  assign data_r[465] = data_r_465_sv2v_reg;
  assign data_r[464] = data_r_464_sv2v_reg;
  assign data_r[463] = data_r_463_sv2v_reg;
  assign data_r[462] = data_r_462_sv2v_reg;
  assign data_r[461] = data_r_461_sv2v_reg;
  assign data_r[460] = data_r_460_sv2v_reg;
  assign data_r[459] = data_r_459_sv2v_reg;
  assign data_r[458] = data_r_458_sv2v_reg;
  assign data_r[457] = data_r_457_sv2v_reg;
  assign data_r[456] = data_r_456_sv2v_reg;
  assign data_r[455] = data_r_455_sv2v_reg;
  assign data_r[454] = data_r_454_sv2v_reg;
  assign data_r[453] = data_r_453_sv2v_reg;
  assign data_r[452] = data_r_452_sv2v_reg;
  assign data_r[451] = data_r_451_sv2v_reg;
  assign data_r[450] = data_r_450_sv2v_reg;
  assign data_r[449] = data_r_449_sv2v_reg;
  assign data_r[448] = data_r_448_sv2v_reg;
  assign data_r[447] = data_r_447_sv2v_reg;
  assign data_r[446] = data_r_446_sv2v_reg;
  assign data_r[445] = data_r_445_sv2v_reg;
  assign data_r[444] = data_r_444_sv2v_reg;
  assign data_r[443] = data_r_443_sv2v_reg;
  assign data_r[442] = data_r_442_sv2v_reg;
  assign data_r[441] = data_r_441_sv2v_reg;
  assign data_r[440] = data_r_440_sv2v_reg;
  assign data_r[439] = data_r_439_sv2v_reg;
  assign data_r[438] = data_r_438_sv2v_reg;
  assign data_r[437] = data_r_437_sv2v_reg;
  assign data_r[436] = data_r_436_sv2v_reg;
  assign data_r[435] = data_r_435_sv2v_reg;
  assign data_r[434] = data_r_434_sv2v_reg;
  assign data_r[433] = data_r_433_sv2v_reg;
  assign data_r[432] = data_r_432_sv2v_reg;
  assign data_r[431] = data_r_431_sv2v_reg;
  assign data_r[430] = data_r_430_sv2v_reg;
  assign data_r[429] = data_r_429_sv2v_reg;
  assign data_r[428] = data_r_428_sv2v_reg;
  assign data_r[427] = data_r_427_sv2v_reg;
  assign data_r[426] = data_r_426_sv2v_reg;
  assign data_r[425] = data_r_425_sv2v_reg;
  assign data_r[424] = data_r_424_sv2v_reg;
  assign data_r[423] = data_r_423_sv2v_reg;
  assign data_r[422] = data_r_422_sv2v_reg;
  assign data_r[421] = data_r_421_sv2v_reg;
  assign data_r[420] = data_r_420_sv2v_reg;
  assign data_r[419] = data_r_419_sv2v_reg;
  assign data_r[418] = data_r_418_sv2v_reg;
  assign data_r[417] = data_r_417_sv2v_reg;
  assign data_r[416] = data_r_416_sv2v_reg;
  assign data_r[415] = data_r_415_sv2v_reg;
  assign data_r[414] = data_r_414_sv2v_reg;
  assign data_r[413] = data_r_413_sv2v_reg;
  assign data_r[412] = data_r_412_sv2v_reg;
  assign data_r[411] = data_r_411_sv2v_reg;
  assign data_r[410] = data_r_410_sv2v_reg;
  assign data_r[409] = data_r_409_sv2v_reg;
  assign data_r[408] = data_r_408_sv2v_reg;
  assign data_r[407] = data_r_407_sv2v_reg;
  assign data_r[406] = data_r_406_sv2v_reg;
  assign data_r[405] = data_r_405_sv2v_reg;
  assign data_r[404] = data_r_404_sv2v_reg;
  assign data_r[403] = data_r_403_sv2v_reg;
  assign data_r[402] = data_r_402_sv2v_reg;
  assign data_r[401] = data_r_401_sv2v_reg;
  assign data_r[400] = data_r_400_sv2v_reg;
  assign data_r[399] = data_r_399_sv2v_reg;
  assign data_r[398] = data_r_398_sv2v_reg;
  assign data_r[397] = data_r_397_sv2v_reg;
  assign data_r[396] = data_r_396_sv2v_reg;
  assign data_r[395] = data_r_395_sv2v_reg;
  assign data_r[394] = data_r_394_sv2v_reg;
  assign data_r[393] = data_r_393_sv2v_reg;
  assign data_r[392] = data_r_392_sv2v_reg;
  assign data_r[391] = data_r_391_sv2v_reg;
  assign data_r[390] = data_r_390_sv2v_reg;
  assign data_r[389] = data_r_389_sv2v_reg;
  assign data_r[388] = data_r_388_sv2v_reg;
  assign data_r[387] = data_r_387_sv2v_reg;
  assign data_r[386] = data_r_386_sv2v_reg;
  assign data_r[385] = data_r_385_sv2v_reg;
  assign data_r[384] = data_r_384_sv2v_reg;
  assign data_r[383] = data_r_383_sv2v_reg;
  assign data_r[382] = data_r_382_sv2v_reg;
  assign data_r[381] = data_r_381_sv2v_reg;
  assign data_r[380] = data_r_380_sv2v_reg;
  assign data_r[379] = data_r_379_sv2v_reg;
  assign data_r[378] = data_r_378_sv2v_reg;
  assign data_r[377] = data_r_377_sv2v_reg;
  assign data_r[376] = data_r_376_sv2v_reg;
  assign data_r[375] = data_r_375_sv2v_reg;
  assign data_r[374] = data_r_374_sv2v_reg;
  assign data_r[373] = data_r_373_sv2v_reg;
  assign data_r[372] = data_r_372_sv2v_reg;
  assign data_r[371] = data_r_371_sv2v_reg;
  assign data_r[370] = data_r_370_sv2v_reg;
  assign data_r[369] = data_r_369_sv2v_reg;
  assign data_r[368] = data_r_368_sv2v_reg;
  assign data_r[367] = data_r_367_sv2v_reg;
  assign data_r[366] = data_r_366_sv2v_reg;
  assign data_r[365] = data_r_365_sv2v_reg;
  assign data_r[364] = data_r_364_sv2v_reg;
  assign data_r[363] = data_r_363_sv2v_reg;
  assign data_r[362] = data_r_362_sv2v_reg;
  assign data_r[361] = data_r_361_sv2v_reg;
  assign data_r[360] = data_r_360_sv2v_reg;
  assign data_r[359] = data_r_359_sv2v_reg;
  assign data_r[358] = data_r_358_sv2v_reg;
  assign data_r[357] = data_r_357_sv2v_reg;
  assign data_r[356] = data_r_356_sv2v_reg;
  assign data_r[355] = data_r_355_sv2v_reg;
  assign data_r[354] = data_r_354_sv2v_reg;
  assign data_r[353] = data_r_353_sv2v_reg;
  assign data_r[352] = data_r_352_sv2v_reg;
  assign data_r[351] = data_r_351_sv2v_reg;
  assign data_r[350] = data_r_350_sv2v_reg;
  assign data_r[349] = data_r_349_sv2v_reg;
  assign data_r[348] = data_r_348_sv2v_reg;
  assign data_r[347] = data_r_347_sv2v_reg;
  assign data_r[346] = data_r_346_sv2v_reg;
  assign data_r[345] = data_r_345_sv2v_reg;
  assign data_r[344] = data_r_344_sv2v_reg;
  assign data_r[343] = data_r_343_sv2v_reg;
  assign data_r[342] = data_r_342_sv2v_reg;
  assign data_r[341] = data_r_341_sv2v_reg;
  assign data_r[340] = data_r_340_sv2v_reg;
  assign data_r[339] = data_r_339_sv2v_reg;
  assign data_r[338] = data_r_338_sv2v_reg;
  assign data_r[337] = data_r_337_sv2v_reg;
  assign data_r[336] = data_r_336_sv2v_reg;
  assign data_r[335] = data_r_335_sv2v_reg;
  assign data_r[334] = data_r_334_sv2v_reg;
  assign data_r[333] = data_r_333_sv2v_reg;
  assign data_r[332] = data_r_332_sv2v_reg;
  assign data_r[331] = data_r_331_sv2v_reg;
  assign data_r[330] = data_r_330_sv2v_reg;
  assign data_r[329] = data_r_329_sv2v_reg;
  assign data_r[328] = data_r_328_sv2v_reg;
  assign data_r[327] = data_r_327_sv2v_reg;
  assign data_r[326] = data_r_326_sv2v_reg;
  assign data_r[325] = data_r_325_sv2v_reg;
  assign data_r[324] = data_r_324_sv2v_reg;
  assign data_r[323] = data_r_323_sv2v_reg;
  assign data_r[322] = data_r_322_sv2v_reg;
  assign data_r[321] = data_r_321_sv2v_reg;
  assign data_r[320] = data_r_320_sv2v_reg;
  assign data_r[319] = data_r_319_sv2v_reg;
  assign data_r[318] = data_r_318_sv2v_reg;
  assign data_r[317] = data_r_317_sv2v_reg;
  assign data_r[316] = data_r_316_sv2v_reg;
  assign data_r[315] = data_r_315_sv2v_reg;
  assign data_r[314] = data_r_314_sv2v_reg;
  assign data_r[313] = data_r_313_sv2v_reg;
  assign data_r[312] = data_r_312_sv2v_reg;
  assign data_r[311] = data_r_311_sv2v_reg;
  assign data_r[310] = data_r_310_sv2v_reg;
  assign data_r[309] = data_r_309_sv2v_reg;
  assign data_r[308] = data_r_308_sv2v_reg;
  assign data_r[307] = data_r_307_sv2v_reg;
  assign data_r[306] = data_r_306_sv2v_reg;
  assign data_r[305] = data_r_305_sv2v_reg;
  assign data_r[304] = data_r_304_sv2v_reg;
  assign data_r[303] = data_r_303_sv2v_reg;
  assign data_r[302] = data_r_302_sv2v_reg;
  assign data_r[301] = data_r_301_sv2v_reg;
  assign data_r[300] = data_r_300_sv2v_reg;
  assign data_r[299] = data_r_299_sv2v_reg;
  assign data_r[298] = data_r_298_sv2v_reg;
  assign data_r[297] = data_r_297_sv2v_reg;
  assign data_r[296] = data_r_296_sv2v_reg;
  assign data_r[295] = data_r_295_sv2v_reg;
  assign data_r[294] = data_r_294_sv2v_reg;
  assign data_r[293] = data_r_293_sv2v_reg;
  assign data_r[292] = data_r_292_sv2v_reg;
  assign data_r[291] = data_r_291_sv2v_reg;
  assign data_r[290] = data_r_290_sv2v_reg;
  assign data_r[289] = data_r_289_sv2v_reg;
  assign data_r[288] = data_r_288_sv2v_reg;
  assign data_r[287] = data_r_287_sv2v_reg;
  assign data_r[286] = data_r_286_sv2v_reg;
  assign data_r[285] = data_r_285_sv2v_reg;
  assign data_r[284] = data_r_284_sv2v_reg;
  assign data_r[283] = data_r_283_sv2v_reg;
  assign data_r[282] = data_r_282_sv2v_reg;
  assign data_r[281] = data_r_281_sv2v_reg;
  assign data_r[280] = data_r_280_sv2v_reg;
  assign data_r[279] = data_r_279_sv2v_reg;
  assign data_r[278] = data_r_278_sv2v_reg;
  assign data_r[277] = data_r_277_sv2v_reg;
  assign data_r[276] = data_r_276_sv2v_reg;
  assign data_r[275] = data_r_275_sv2v_reg;
  assign data_r[274] = data_r_274_sv2v_reg;
  assign data_r[273] = data_r_273_sv2v_reg;
  assign data_r[272] = data_r_272_sv2v_reg;
  assign data_r[271] = data_r_271_sv2v_reg;
  assign data_r[270] = data_r_270_sv2v_reg;
  assign data_r[269] = data_r_269_sv2v_reg;
  assign data_r[268] = data_r_268_sv2v_reg;
  assign data_r[267] = data_r_267_sv2v_reg;
  assign data_r[266] = data_r_266_sv2v_reg;
  assign data_r[265] = data_r_265_sv2v_reg;
  assign data_r[264] = data_r_264_sv2v_reg;
  assign data_r[263] = data_r_263_sv2v_reg;
  assign data_r[262] = data_r_262_sv2v_reg;
  assign data_r[261] = data_r_261_sv2v_reg;
  assign data_r[260] = data_r_260_sv2v_reg;
  assign data_r[259] = data_r_259_sv2v_reg;
  assign data_r[258] = data_r_258_sv2v_reg;
  assign data_r[257] = data_r_257_sv2v_reg;
  assign data_r[256] = data_r_256_sv2v_reg;
  assign data_r[255] = data_r_255_sv2v_reg;
  assign data_r[254] = data_r_254_sv2v_reg;
  assign data_r[253] = data_r_253_sv2v_reg;
  assign data_r[252] = data_r_252_sv2v_reg;
  assign data_r[251] = data_r_251_sv2v_reg;
  assign data_r[250] = data_r_250_sv2v_reg;
  assign data_r[249] = data_r_249_sv2v_reg;
  assign data_r[248] = data_r_248_sv2v_reg;
  assign data_r[247] = data_r_247_sv2v_reg;
  assign data_r[246] = data_r_246_sv2v_reg;
  assign data_r[245] = data_r_245_sv2v_reg;
  assign data_r[244] = data_r_244_sv2v_reg;
  assign data_r[243] = data_r_243_sv2v_reg;
  assign data_r[242] = data_r_242_sv2v_reg;
  assign data_r[241] = data_r_241_sv2v_reg;
  assign data_r[240] = data_r_240_sv2v_reg;
  assign data_r[239] = data_r_239_sv2v_reg;
  assign data_r[238] = data_r_238_sv2v_reg;
  assign data_r[237] = data_r_237_sv2v_reg;
  assign data_r[236] = data_r_236_sv2v_reg;
  assign data_r[235] = data_r_235_sv2v_reg;
  assign data_r[234] = data_r_234_sv2v_reg;
  assign data_r[233] = data_r_233_sv2v_reg;
  assign data_r[232] = data_r_232_sv2v_reg;
  assign data_r[231] = data_r_231_sv2v_reg;
  assign data_r[230] = data_r_230_sv2v_reg;
  assign data_r[229] = data_r_229_sv2v_reg;
  assign data_r[228] = data_r_228_sv2v_reg;
  assign data_r[227] = data_r_227_sv2v_reg;
  assign data_r[226] = data_r_226_sv2v_reg;
  assign data_r[225] = data_r_225_sv2v_reg;
  assign data_r[224] = data_r_224_sv2v_reg;
  assign data_r[223] = data_r_223_sv2v_reg;
  assign data_r[222] = data_r_222_sv2v_reg;
  assign data_r[221] = data_r_221_sv2v_reg;
  assign data_r[220] = data_r_220_sv2v_reg;
  assign data_r[219] = data_r_219_sv2v_reg;
  assign data_r[218] = data_r_218_sv2v_reg;
  assign data_r[217] = data_r_217_sv2v_reg;
  assign data_r[216] = data_r_216_sv2v_reg;
  assign data_r[215] = data_r_215_sv2v_reg;
  assign data_r[214] = data_r_214_sv2v_reg;
  assign data_r[213] = data_r_213_sv2v_reg;
  assign data_r[212] = data_r_212_sv2v_reg;
  assign data_r[211] = data_r_211_sv2v_reg;
  assign data_r[210] = data_r_210_sv2v_reg;
  assign data_r[209] = data_r_209_sv2v_reg;
  assign data_r[208] = data_r_208_sv2v_reg;
  assign data_r[207] = data_r_207_sv2v_reg;
  assign data_r[206] = data_r_206_sv2v_reg;
  assign data_r[205] = data_r_205_sv2v_reg;
  assign data_r[204] = data_r_204_sv2v_reg;
  assign data_r[203] = data_r_203_sv2v_reg;
  assign data_r[202] = data_r_202_sv2v_reg;
  assign data_r[201] = data_r_201_sv2v_reg;
  assign data_r[200] = data_r_200_sv2v_reg;
  assign data_r[199] = data_r_199_sv2v_reg;
  assign data_r[198] = data_r_198_sv2v_reg;
  assign data_r[197] = data_r_197_sv2v_reg;
  assign data_r[196] = data_r_196_sv2v_reg;
  assign data_r[195] = data_r_195_sv2v_reg;
  assign data_r[194] = data_r_194_sv2v_reg;
  assign data_r[193] = data_r_193_sv2v_reg;
  assign data_r[192] = data_r_192_sv2v_reg;
  assign data_r[191] = data_r_191_sv2v_reg;
  assign data_r[190] = data_r_190_sv2v_reg;
  assign data_r[189] = data_r_189_sv2v_reg;
  assign data_r[188] = data_r_188_sv2v_reg;
  assign data_r[187] = data_r_187_sv2v_reg;
  assign data_r[186] = data_r_186_sv2v_reg;
  assign data_r[185] = data_r_185_sv2v_reg;
  assign data_r[184] = data_r_184_sv2v_reg;
  assign data_r[183] = data_r_183_sv2v_reg;
  assign data_r[182] = data_r_182_sv2v_reg;
  assign data_r[181] = data_r_181_sv2v_reg;
  assign data_r[180] = data_r_180_sv2v_reg;
  assign data_r[179] = data_r_179_sv2v_reg;
  assign data_r[178] = data_r_178_sv2v_reg;
  assign data_r[177] = data_r_177_sv2v_reg;
  assign data_r[176] = data_r_176_sv2v_reg;
  assign data_r[175] = data_r_175_sv2v_reg;
  assign data_r[174] = data_r_174_sv2v_reg;
  assign data_r[173] = data_r_173_sv2v_reg;
  assign data_r[172] = data_r_172_sv2v_reg;
  assign data_r[171] = data_r_171_sv2v_reg;
  assign data_r[170] = data_r_170_sv2v_reg;
  assign data_r[169] = data_r_169_sv2v_reg;
  assign data_r[168] = data_r_168_sv2v_reg;
  assign data_r[167] = data_r_167_sv2v_reg;
  assign data_r[166] = data_r_166_sv2v_reg;
  assign data_r[165] = data_r_165_sv2v_reg;
  assign data_r[164] = data_r_164_sv2v_reg;
  assign data_r[163] = data_r_163_sv2v_reg;
  assign data_r[162] = data_r_162_sv2v_reg;
  assign data_r[161] = data_r_161_sv2v_reg;
  assign data_r[160] = data_r_160_sv2v_reg;
  assign data_r[159] = data_r_159_sv2v_reg;
  assign data_r[158] = data_r_158_sv2v_reg;
  assign data_r[157] = data_r_157_sv2v_reg;
  assign data_r[156] = data_r_156_sv2v_reg;
  assign data_r[155] = data_r_155_sv2v_reg;
  assign data_r[154] = data_r_154_sv2v_reg;
  assign data_r[153] = data_r_153_sv2v_reg;
  assign data_r[152] = data_r_152_sv2v_reg;
  assign data_r[151] = data_r_151_sv2v_reg;
  assign data_r[150] = data_r_150_sv2v_reg;
  assign data_r[149] = data_r_149_sv2v_reg;
  assign data_r[148] = data_r_148_sv2v_reg;
  assign data_r[147] = data_r_147_sv2v_reg;
  assign data_r[146] = data_r_146_sv2v_reg;
  assign data_r[145] = data_r_145_sv2v_reg;
  assign data_r[144] = data_r_144_sv2v_reg;
  assign data_r[143] = data_r_143_sv2v_reg;
  assign data_r[142] = data_r_142_sv2v_reg;
  assign data_r[141] = data_r_141_sv2v_reg;
  assign data_r[140] = data_r_140_sv2v_reg;
  assign data_r[139] = data_r_139_sv2v_reg;
  assign data_r[138] = data_r_138_sv2v_reg;
  assign data_r[137] = data_r_137_sv2v_reg;
  assign data_r[136] = data_r_136_sv2v_reg;
  assign data_r[135] = data_r_135_sv2v_reg;
  assign data_r[134] = data_r_134_sv2v_reg;
  assign data_r[133] = data_r_133_sv2v_reg;
  assign data_r[132] = data_r_132_sv2v_reg;
  assign data_r[131] = data_r_131_sv2v_reg;
  assign data_r[130] = data_r_130_sv2v_reg;
  assign data_r[129] = data_r_129_sv2v_reg;
  assign data_r[128] = data_r_128_sv2v_reg;
  assign data_r[127] = data_r_127_sv2v_reg;
  assign data_r[126] = data_r_126_sv2v_reg;
  assign data_r[125] = data_r_125_sv2v_reg;
  assign data_r[124] = data_r_124_sv2v_reg;
  assign data_r[123] = data_r_123_sv2v_reg;
  assign data_r[122] = data_r_122_sv2v_reg;
  assign data_r[121] = data_r_121_sv2v_reg;
  assign data_r[120] = data_r_120_sv2v_reg;
  assign data_r[119] = data_r_119_sv2v_reg;
  assign data_r[118] = data_r_118_sv2v_reg;
  assign data_r[117] = data_r_117_sv2v_reg;
  assign data_r[116] = data_r_116_sv2v_reg;
  assign data_r[115] = data_r_115_sv2v_reg;
  assign data_r[114] = data_r_114_sv2v_reg;
  assign data_r[113] = data_r_113_sv2v_reg;
  assign data_r[112] = data_r_112_sv2v_reg;
  assign data_r[111] = data_r_111_sv2v_reg;
  assign data_r[110] = data_r_110_sv2v_reg;
  assign data_r[109] = data_r_109_sv2v_reg;
  assign data_r[108] = data_r_108_sv2v_reg;
  assign data_r[107] = data_r_107_sv2v_reg;
  assign data_r[106] = data_r_106_sv2v_reg;
  assign data_r[105] = data_r_105_sv2v_reg;
  assign data_r[104] = data_r_104_sv2v_reg;
  assign data_r[103] = data_r_103_sv2v_reg;
  assign data_r[102] = data_r_102_sv2v_reg;
  assign data_r[101] = data_r_101_sv2v_reg;
  assign data_r[100] = data_r_100_sv2v_reg;
  assign data_r[99] = data_r_99_sv2v_reg;
  assign data_r[98] = data_r_98_sv2v_reg;
  assign data_r[97] = data_r_97_sv2v_reg;
  assign data_r[96] = data_r_96_sv2v_reg;
  assign data_r[95] = data_r_95_sv2v_reg;
  assign data_r[94] = data_r_94_sv2v_reg;
  assign data_r[93] = data_r_93_sv2v_reg;
  assign data_r[92] = data_r_92_sv2v_reg;
  assign data_r[91] = data_r_91_sv2v_reg;
  assign data_r[90] = data_r_90_sv2v_reg;
  assign data_r[89] = data_r_89_sv2v_reg;
  assign data_r[88] = data_r_88_sv2v_reg;
  assign data_r[87] = data_r_87_sv2v_reg;
  assign data_r[86] = data_r_86_sv2v_reg;
  assign data_r[85] = data_r_85_sv2v_reg;
  assign data_r[84] = data_r_84_sv2v_reg;
  assign data_r[83] = data_r_83_sv2v_reg;
  assign data_r[82] = data_r_82_sv2v_reg;
  assign data_r[81] = data_r_81_sv2v_reg;
  assign data_r[80] = data_r_80_sv2v_reg;
  assign data_r[79] = data_r_79_sv2v_reg;
  assign data_r[78] = data_r_78_sv2v_reg;
  assign data_r[77] = data_r_77_sv2v_reg;
  assign data_r[76] = data_r_76_sv2v_reg;
  assign data_r[75] = data_r_75_sv2v_reg;
  assign data_r[74] = data_r_74_sv2v_reg;
  assign data_r[73] = data_r_73_sv2v_reg;
  assign data_r[72] = data_r_72_sv2v_reg;
  assign data_r[71] = data_r_71_sv2v_reg;
  assign data_r[70] = data_r_70_sv2v_reg;
  assign data_r[69] = data_r_69_sv2v_reg;
  assign data_r[68] = data_r_68_sv2v_reg;
  assign data_r[67] = data_r_67_sv2v_reg;
  assign data_r[66] = data_r_66_sv2v_reg;
  assign data_r[65] = data_r_65_sv2v_reg;
  assign data_r[64] = data_r_64_sv2v_reg;
  assign data_r[63] = data_r_63_sv2v_reg;
  assign data_r[62] = data_r_62_sv2v_reg;
  assign data_r[61] = data_r_61_sv2v_reg;
  assign data_r[60] = data_r_60_sv2v_reg;
  assign data_r[59] = data_r_59_sv2v_reg;
  assign data_r[58] = data_r_58_sv2v_reg;
  assign data_r[57] = data_r_57_sv2v_reg;
  assign data_r[56] = data_r_56_sv2v_reg;
  assign data_r[55] = data_r_55_sv2v_reg;
  assign data_r[54] = data_r_54_sv2v_reg;
  assign data_r[53] = data_r_53_sv2v_reg;
  assign data_r[52] = data_r_52_sv2v_reg;
  assign data_r[51] = data_r_51_sv2v_reg;
  assign data_r[50] = data_r_50_sv2v_reg;
  assign data_r[49] = data_r_49_sv2v_reg;
  assign data_r[48] = data_r_48_sv2v_reg;
  assign data_r[47] = data_r_47_sv2v_reg;
  assign data_r[46] = data_r_46_sv2v_reg;
  assign data_r[45] = data_r_45_sv2v_reg;
  assign data_r[44] = data_r_44_sv2v_reg;
  assign data_r[43] = data_r_43_sv2v_reg;
  assign data_r[42] = data_r_42_sv2v_reg;
  assign data_r[41] = data_r_41_sv2v_reg;
  assign data_r[40] = data_r_40_sv2v_reg;
  assign data_r[39] = data_r_39_sv2v_reg;
  assign data_r[38] = data_r_38_sv2v_reg;
  assign data_r[37] = data_r_37_sv2v_reg;
  assign data_r[36] = data_r_36_sv2v_reg;
  assign data_r[35] = data_r_35_sv2v_reg;
  assign data_r[34] = data_r_34_sv2v_reg;
  assign data_r[33] = data_r_33_sv2v_reg;
  assign data_r[32] = data_r_32_sv2v_reg;
  assign data_r[31] = data_r_31_sv2v_reg;
  assign data_r[30] = data_r_30_sv2v_reg;
  assign data_r[29] = data_r_29_sv2v_reg;
  assign data_r[28] = data_r_28_sv2v_reg;
  assign data_r[27] = data_r_27_sv2v_reg;
  assign data_r[26] = data_r_26_sv2v_reg;
  assign data_r[25] = data_r_25_sv2v_reg;
  assign data_r[24] = data_r_24_sv2v_reg;
  assign data_r[23] = data_r_23_sv2v_reg;
  assign data_r[22] = data_r_22_sv2v_reg;
  assign data_r[21] = data_r_21_sv2v_reg;
  assign data_r[20] = data_r_20_sv2v_reg;
  assign data_r[19] = data_r_19_sv2v_reg;
  assign data_r[18] = data_r_18_sv2v_reg;
  assign data_r[17] = data_r_17_sv2v_reg;
  assign data_r[16] = data_r_16_sv2v_reg;
  assign data_r[15] = data_r_15_sv2v_reg;
  assign data_r[14] = data_r_14_sv2v_reg;
  assign data_r[13] = data_r_13_sv2v_reg;
  assign data_r[12] = data_r_12_sv2v_reg;
  assign data_r[11] = data_r_11_sv2v_reg;
  assign data_r[10] = data_r_10_sv2v_reg;
  assign data_r[9] = data_r_9_sv2v_reg;
  assign data_r[8] = data_r_8_sv2v_reg;
  assign data_r[7] = data_r_7_sv2v_reg;
  assign data_r[6] = data_r_6_sv2v_reg;
  assign data_r[5] = data_r_5_sv2v_reg;
  assign data_r[4] = data_r_4_sv2v_reg;
  assign data_r[3] = data_r_3_sv2v_reg;
  assign data_r[2] = data_r_2_sv2v_reg;
  assign data_r[1] = data_r_1_sv2v_reg;
  assign data_r[0] = data_r_0_sv2v_reg;
  assign data_nn[15] = (N732)? data_o[15] : 
                       (N734)? data_o[31] : 
                       (N736)? data_o[47] : 
                       (N738)? data_o[63] : 
                       (N740)? data_o[79] : 
                       (N742)? data_o[95] : 
                       (N744)? data_o[111] : 
                       (N746)? data_o[127] : 
                       (N748)? data_o[143] : 
                       (N750)? data_o[159] : 
                       (N752)? data_o[175] : 
                       (N754)? data_o[191] : 
                       (N756)? data_o[207] : 
                       (N758)? data_o[223] : 
                       (N760)? data_o[239] : 
                       (N762)? data_o[255] : 
                       (N764)? data_o[271] : 
                       (N766)? data_o[287] : 
                       (N768)? data_o[303] : 
                       (N770)? data_o[319] : 
                       (N772)? data_o[335] : 
                       (N774)? data_o[351] : 
                       (N776)? data_o[367] : 
                       (N778)? data_o[383] : 
                       (N780)? data_o[399] : 
                       (N782)? data_o[415] : 
                       (N784)? data_o[431] : 
                       (N786)? data_o[447] : 
                       (N788)? data_o[463] : 
                       (N790)? data_o[479] : 
                       (N792)? data_o[495] : 
                       (N794)? data_o[511] : 
                       (N733)? data_n_32__15_ : 
                       (N735)? data_n_33__15_ : 
                       (N737)? data_n_34__15_ : 
                       (N739)? data_n_35__15_ : 
                       (N741)? data_n_36__15_ : 
                       (N743)? data_n_37__15_ : 
                       (N745)? data_n_38__15_ : 
                       (N747)? data_n_39__15_ : 
                       (N749)? data_n_40__15_ : 
                       (N751)? data_n_41__15_ : 
                       (N753)? data_n_42__15_ : 
                       (N755)? data_n_43__15_ : 
                       (N757)? data_n_44__15_ : 
                       (N759)? data_n_45__15_ : 
                       (N761)? data_n_46__15_ : 
                       (N763)? data_n_47__15_ : 
                       (N765)? data_n_48__15_ : 
                       (N767)? data_n_49__15_ : 
                       (N769)? data_n_50__15_ : 
                       (N771)? data_n_51__15_ : 
                       (N773)? data_n_52__15_ : 
                       (N775)? data_n_53__15_ : 
                       (N777)? data_n_54__15_ : 
                       (N779)? data_n_55__15_ : 
                       (N781)? data_n_56__15_ : 
                       (N783)? data_n_57__15_ : 
                       (N785)? data_n_58__15_ : 
                       (N787)? data_n_59__15_ : 
                       (N789)? data_n_60__15_ : 
                       (N791)? data_n_61__15_ : 
                       (N793)? data_n_62__15_ : 
                       (N795)? data_n_63__15_ : 1'b0;
  assign data_nn[14] = (N732)? data_o[14] : 
                       (N734)? data_o[30] : 
                       (N736)? data_o[46] : 
                       (N738)? data_o[62] : 
                       (N740)? data_o[78] : 
                       (N742)? data_o[94] : 
                       (N744)? data_o[110] : 
                       (N746)? data_o[126] : 
                       (N748)? data_o[142] : 
                       (N750)? data_o[158] : 
                       (N752)? data_o[174] : 
                       (N754)? data_o[190] : 
                       (N756)? data_o[206] : 
                       (N758)? data_o[222] : 
                       (N760)? data_o[238] : 
                       (N762)? data_o[254] : 
                       (N764)? data_o[270] : 
                       (N766)? data_o[286] : 
                       (N768)? data_o[302] : 
                       (N770)? data_o[318] : 
                       (N772)? data_o[334] : 
                       (N774)? data_o[350] : 
                       (N776)? data_o[366] : 
                       (N778)? data_o[382] : 
                       (N780)? data_o[398] : 
                       (N782)? data_o[414] : 
                       (N784)? data_o[430] : 
                       (N786)? data_o[446] : 
                       (N788)? data_o[462] : 
                       (N790)? data_o[478] : 
                       (N792)? data_o[494] : 
                       (N794)? data_o[510] : 
                       (N733)? data_n_32__14_ : 
                       (N735)? data_n_33__14_ : 
                       (N737)? data_n_34__14_ : 
                       (N739)? data_n_35__14_ : 
                       (N741)? data_n_36__14_ : 
                       (N743)? data_n_37__14_ : 
                       (N745)? data_n_38__14_ : 
                       (N747)? data_n_39__14_ : 
                       (N749)? data_n_40__14_ : 
                       (N751)? data_n_41__14_ : 
                       (N753)? data_n_42__14_ : 
                       (N755)? data_n_43__14_ : 
                       (N757)? data_n_44__14_ : 
                       (N759)? data_n_45__14_ : 
                       (N761)? data_n_46__14_ : 
                       (N763)? data_n_47__14_ : 
                       (N765)? data_n_48__14_ : 
                       (N767)? data_n_49__14_ : 
                       (N769)? data_n_50__14_ : 
                       (N771)? data_n_51__14_ : 
                       (N773)? data_n_52__14_ : 
                       (N775)? data_n_53__14_ : 
                       (N777)? data_n_54__14_ : 
                       (N779)? data_n_55__14_ : 
                       (N781)? data_n_56__14_ : 
                       (N783)? data_n_57__14_ : 
                       (N785)? data_n_58__14_ : 
                       (N787)? data_n_59__14_ : 
                       (N789)? data_n_60__14_ : 
                       (N791)? data_n_61__14_ : 
                       (N793)? data_n_62__14_ : 
                       (N795)? data_n_63__14_ : 1'b0;
  assign data_nn[13] = (N732)? data_o[13] : 
                       (N734)? data_o[29] : 
                       (N736)? data_o[45] : 
                       (N738)? data_o[61] : 
                       (N740)? data_o[77] : 
                       (N742)? data_o[93] : 
                       (N744)? data_o[109] : 
                       (N746)? data_o[125] : 
                       (N748)? data_o[141] : 
                       (N750)? data_o[157] : 
                       (N752)? data_o[173] : 
                       (N754)? data_o[189] : 
                       (N756)? data_o[205] : 
                       (N758)? data_o[221] : 
                       (N760)? data_o[237] : 
                       (N762)? data_o[253] : 
                       (N764)? data_o[269] : 
                       (N766)? data_o[285] : 
                       (N768)? data_o[301] : 
                       (N770)? data_o[317] : 
                       (N772)? data_o[333] : 
                       (N774)? data_o[349] : 
                       (N776)? data_o[365] : 
                       (N778)? data_o[381] : 
                       (N780)? data_o[397] : 
                       (N782)? data_o[413] : 
                       (N784)? data_o[429] : 
                       (N786)? data_o[445] : 
                       (N788)? data_o[461] : 
                       (N790)? data_o[477] : 
                       (N792)? data_o[493] : 
                       (N794)? data_o[509] : 
                       (N733)? data_n_32__13_ : 
                       (N735)? data_n_33__13_ : 
                       (N737)? data_n_34__13_ : 
                       (N739)? data_n_35__13_ : 
                       (N741)? data_n_36__13_ : 
                       (N743)? data_n_37__13_ : 
                       (N745)? data_n_38__13_ : 
                       (N747)? data_n_39__13_ : 
                       (N749)? data_n_40__13_ : 
                       (N751)? data_n_41__13_ : 
                       (N753)? data_n_42__13_ : 
                       (N755)? data_n_43__13_ : 
                       (N757)? data_n_44__13_ : 
                       (N759)? data_n_45__13_ : 
                       (N761)? data_n_46__13_ : 
                       (N763)? data_n_47__13_ : 
                       (N765)? data_n_48__13_ : 
                       (N767)? data_n_49__13_ : 
                       (N769)? data_n_50__13_ : 
                       (N771)? data_n_51__13_ : 
                       (N773)? data_n_52__13_ : 
                       (N775)? data_n_53__13_ : 
                       (N777)? data_n_54__13_ : 
                       (N779)? data_n_55__13_ : 
                       (N781)? data_n_56__13_ : 
                       (N783)? data_n_57__13_ : 
                       (N785)? data_n_58__13_ : 
                       (N787)? data_n_59__13_ : 
                       (N789)? data_n_60__13_ : 
                       (N791)? data_n_61__13_ : 
                       (N793)? data_n_62__13_ : 
                       (N795)? data_n_63__13_ : 1'b0;
  assign data_nn[12] = (N732)? data_o[12] : 
                       (N734)? data_o[28] : 
                       (N736)? data_o[44] : 
                       (N738)? data_o[60] : 
                       (N740)? data_o[76] : 
                       (N742)? data_o[92] : 
                       (N744)? data_o[108] : 
                       (N746)? data_o[124] : 
                       (N748)? data_o[140] : 
                       (N750)? data_o[156] : 
                       (N752)? data_o[172] : 
                       (N754)? data_o[188] : 
                       (N756)? data_o[204] : 
                       (N758)? data_o[220] : 
                       (N760)? data_o[236] : 
                       (N762)? data_o[252] : 
                       (N764)? data_o[268] : 
                       (N766)? data_o[284] : 
                       (N768)? data_o[300] : 
                       (N770)? data_o[316] : 
                       (N772)? data_o[332] : 
                       (N774)? data_o[348] : 
                       (N776)? data_o[364] : 
                       (N778)? data_o[380] : 
                       (N780)? data_o[396] : 
                       (N782)? data_o[412] : 
                       (N784)? data_o[428] : 
                       (N786)? data_o[444] : 
                       (N788)? data_o[460] : 
                       (N790)? data_o[476] : 
                       (N792)? data_o[492] : 
                       (N794)? data_o[508] : 
                       (N733)? data_n_32__12_ : 
                       (N735)? data_n_33__12_ : 
                       (N737)? data_n_34__12_ : 
                       (N739)? data_n_35__12_ : 
                       (N741)? data_n_36__12_ : 
                       (N743)? data_n_37__12_ : 
                       (N745)? data_n_38__12_ : 
                       (N747)? data_n_39__12_ : 
                       (N749)? data_n_40__12_ : 
                       (N751)? data_n_41__12_ : 
                       (N753)? data_n_42__12_ : 
                       (N755)? data_n_43__12_ : 
                       (N757)? data_n_44__12_ : 
                       (N759)? data_n_45__12_ : 
                       (N761)? data_n_46__12_ : 
                       (N763)? data_n_47__12_ : 
                       (N765)? data_n_48__12_ : 
                       (N767)? data_n_49__12_ : 
                       (N769)? data_n_50__12_ : 
                       (N771)? data_n_51__12_ : 
                       (N773)? data_n_52__12_ : 
                       (N775)? data_n_53__12_ : 
                       (N777)? data_n_54__12_ : 
                       (N779)? data_n_55__12_ : 
                       (N781)? data_n_56__12_ : 
                       (N783)? data_n_57__12_ : 
                       (N785)? data_n_58__12_ : 
                       (N787)? data_n_59__12_ : 
                       (N789)? data_n_60__12_ : 
                       (N791)? data_n_61__12_ : 
                       (N793)? data_n_62__12_ : 
                       (N795)? data_n_63__12_ : 1'b0;
  assign data_nn[11] = (N732)? data_o[11] : 
                       (N734)? data_o[27] : 
                       (N736)? data_o[43] : 
                       (N738)? data_o[59] : 
                       (N740)? data_o[75] : 
                       (N742)? data_o[91] : 
                       (N744)? data_o[107] : 
                       (N746)? data_o[123] : 
                       (N748)? data_o[139] : 
                       (N750)? data_o[155] : 
                       (N752)? data_o[171] : 
                       (N754)? data_o[187] : 
                       (N756)? data_o[203] : 
                       (N758)? data_o[219] : 
                       (N760)? data_o[235] : 
                       (N762)? data_o[251] : 
                       (N764)? data_o[267] : 
                       (N766)? data_o[283] : 
                       (N768)? data_o[299] : 
                       (N770)? data_o[315] : 
                       (N772)? data_o[331] : 
                       (N774)? data_o[347] : 
                       (N776)? data_o[363] : 
                       (N778)? data_o[379] : 
                       (N780)? data_o[395] : 
                       (N782)? data_o[411] : 
                       (N784)? data_o[427] : 
                       (N786)? data_o[443] : 
                       (N788)? data_o[459] : 
                       (N790)? data_o[475] : 
                       (N792)? data_o[491] : 
                       (N794)? data_o[507] : 
                       (N733)? data_n_32__11_ : 
                       (N735)? data_n_33__11_ : 
                       (N737)? data_n_34__11_ : 
                       (N739)? data_n_35__11_ : 
                       (N741)? data_n_36__11_ : 
                       (N743)? data_n_37__11_ : 
                       (N745)? data_n_38__11_ : 
                       (N747)? data_n_39__11_ : 
                       (N749)? data_n_40__11_ : 
                       (N751)? data_n_41__11_ : 
                       (N753)? data_n_42__11_ : 
                       (N755)? data_n_43__11_ : 
                       (N757)? data_n_44__11_ : 
                       (N759)? data_n_45__11_ : 
                       (N761)? data_n_46__11_ : 
                       (N763)? data_n_47__11_ : 
                       (N765)? data_n_48__11_ : 
                       (N767)? data_n_49__11_ : 
                       (N769)? data_n_50__11_ : 
                       (N771)? data_n_51__11_ : 
                       (N773)? data_n_52__11_ : 
                       (N775)? data_n_53__11_ : 
                       (N777)? data_n_54__11_ : 
                       (N779)? data_n_55__11_ : 
                       (N781)? data_n_56__11_ : 
                       (N783)? data_n_57__11_ : 
                       (N785)? data_n_58__11_ : 
                       (N787)? data_n_59__11_ : 
                       (N789)? data_n_60__11_ : 
                       (N791)? data_n_61__11_ : 
                       (N793)? data_n_62__11_ : 
                       (N795)? data_n_63__11_ : 1'b0;
  assign data_nn[10] = (N732)? data_o[10] : 
                       (N734)? data_o[26] : 
                       (N736)? data_o[42] : 
                       (N738)? data_o[58] : 
                       (N740)? data_o[74] : 
                       (N742)? data_o[90] : 
                       (N744)? data_o[106] : 
                       (N746)? data_o[122] : 
                       (N748)? data_o[138] : 
                       (N750)? data_o[154] : 
                       (N752)? data_o[170] : 
                       (N754)? data_o[186] : 
                       (N756)? data_o[202] : 
                       (N758)? data_o[218] : 
                       (N760)? data_o[234] : 
                       (N762)? data_o[250] : 
                       (N764)? data_o[266] : 
                       (N766)? data_o[282] : 
                       (N768)? data_o[298] : 
                       (N770)? data_o[314] : 
                       (N772)? data_o[330] : 
                       (N774)? data_o[346] : 
                       (N776)? data_o[362] : 
                       (N778)? data_o[378] : 
                       (N780)? data_o[394] : 
                       (N782)? data_o[410] : 
                       (N784)? data_o[426] : 
                       (N786)? data_o[442] : 
                       (N788)? data_o[458] : 
                       (N790)? data_o[474] : 
                       (N792)? data_o[490] : 
                       (N794)? data_o[506] : 
                       (N733)? data_n_32__10_ : 
                       (N735)? data_n_33__10_ : 
                       (N737)? data_n_34__10_ : 
                       (N739)? data_n_35__10_ : 
                       (N741)? data_n_36__10_ : 
                       (N743)? data_n_37__10_ : 
                       (N745)? data_n_38__10_ : 
                       (N747)? data_n_39__10_ : 
                       (N749)? data_n_40__10_ : 
                       (N751)? data_n_41__10_ : 
                       (N753)? data_n_42__10_ : 
                       (N755)? data_n_43__10_ : 
                       (N757)? data_n_44__10_ : 
                       (N759)? data_n_45__10_ : 
                       (N761)? data_n_46__10_ : 
                       (N763)? data_n_47__10_ : 
                       (N765)? data_n_48__10_ : 
                       (N767)? data_n_49__10_ : 
                       (N769)? data_n_50__10_ : 
                       (N771)? data_n_51__10_ : 
                       (N773)? data_n_52__10_ : 
                       (N775)? data_n_53__10_ : 
                       (N777)? data_n_54__10_ : 
                       (N779)? data_n_55__10_ : 
                       (N781)? data_n_56__10_ : 
                       (N783)? data_n_57__10_ : 
                       (N785)? data_n_58__10_ : 
                       (N787)? data_n_59__10_ : 
                       (N789)? data_n_60__10_ : 
                       (N791)? data_n_61__10_ : 
                       (N793)? data_n_62__10_ : 
                       (N795)? data_n_63__10_ : 1'b0;
  assign data_nn[9] = (N732)? data_o[9] : 
                      (N734)? data_o[25] : 
                      (N736)? data_o[41] : 
                      (N738)? data_o[57] : 
                      (N740)? data_o[73] : 
                      (N742)? data_o[89] : 
                      (N744)? data_o[105] : 
                      (N746)? data_o[121] : 
                      (N748)? data_o[137] : 
                      (N750)? data_o[153] : 
                      (N752)? data_o[169] : 
                      (N754)? data_o[185] : 
                      (N756)? data_o[201] : 
                      (N758)? data_o[217] : 
                      (N760)? data_o[233] : 
                      (N762)? data_o[249] : 
                      (N764)? data_o[265] : 
                      (N766)? data_o[281] : 
                      (N768)? data_o[297] : 
                      (N770)? data_o[313] : 
                      (N772)? data_o[329] : 
                      (N774)? data_o[345] : 
                      (N776)? data_o[361] : 
                      (N778)? data_o[377] : 
                      (N780)? data_o[393] : 
                      (N782)? data_o[409] : 
                      (N784)? data_o[425] : 
                      (N786)? data_o[441] : 
                      (N788)? data_o[457] : 
                      (N790)? data_o[473] : 
                      (N792)? data_o[489] : 
                      (N794)? data_o[505] : 
                      (N733)? data_n_32__9_ : 
                      (N735)? data_n_33__9_ : 
                      (N737)? data_n_34__9_ : 
                      (N739)? data_n_35__9_ : 
                      (N741)? data_n_36__9_ : 
                      (N743)? data_n_37__9_ : 
                      (N745)? data_n_38__9_ : 
                      (N747)? data_n_39__9_ : 
                      (N749)? data_n_40__9_ : 
                      (N751)? data_n_41__9_ : 
                      (N753)? data_n_42__9_ : 
                      (N755)? data_n_43__9_ : 
                      (N757)? data_n_44__9_ : 
                      (N759)? data_n_45__9_ : 
                      (N761)? data_n_46__9_ : 
                      (N763)? data_n_47__9_ : 
                      (N765)? data_n_48__9_ : 
                      (N767)? data_n_49__9_ : 
                      (N769)? data_n_50__9_ : 
                      (N771)? data_n_51__9_ : 
                      (N773)? data_n_52__9_ : 
                      (N775)? data_n_53__9_ : 
                      (N777)? data_n_54__9_ : 
                      (N779)? data_n_55__9_ : 
                      (N781)? data_n_56__9_ : 
                      (N783)? data_n_57__9_ : 
                      (N785)? data_n_58__9_ : 
                      (N787)? data_n_59__9_ : 
                      (N789)? data_n_60__9_ : 
                      (N791)? data_n_61__9_ : 
                      (N793)? data_n_62__9_ : 
                      (N795)? data_n_63__9_ : 1'b0;
  assign data_nn[8] = (N732)? data_o[8] : 
                      (N734)? data_o[24] : 
                      (N736)? data_o[40] : 
                      (N738)? data_o[56] : 
                      (N740)? data_o[72] : 
                      (N742)? data_o[88] : 
                      (N744)? data_o[104] : 
                      (N746)? data_o[120] : 
                      (N748)? data_o[136] : 
                      (N750)? data_o[152] : 
                      (N752)? data_o[168] : 
                      (N754)? data_o[184] : 
                      (N756)? data_o[200] : 
                      (N758)? data_o[216] : 
                      (N760)? data_o[232] : 
                      (N762)? data_o[248] : 
                      (N764)? data_o[264] : 
                      (N766)? data_o[280] : 
                      (N768)? data_o[296] : 
                      (N770)? data_o[312] : 
                      (N772)? data_o[328] : 
                      (N774)? data_o[344] : 
                      (N776)? data_o[360] : 
                      (N778)? data_o[376] : 
                      (N780)? data_o[392] : 
                      (N782)? data_o[408] : 
                      (N784)? data_o[424] : 
                      (N786)? data_o[440] : 
                      (N788)? data_o[456] : 
                      (N790)? data_o[472] : 
                      (N792)? data_o[488] : 
                      (N794)? data_o[504] : 
                      (N733)? data_n_32__8_ : 
                      (N735)? data_n_33__8_ : 
                      (N737)? data_n_34__8_ : 
                      (N739)? data_n_35__8_ : 
                      (N741)? data_n_36__8_ : 
                      (N743)? data_n_37__8_ : 
                      (N745)? data_n_38__8_ : 
                      (N747)? data_n_39__8_ : 
                      (N749)? data_n_40__8_ : 
                      (N751)? data_n_41__8_ : 
                      (N753)? data_n_42__8_ : 
                      (N755)? data_n_43__8_ : 
                      (N757)? data_n_44__8_ : 
                      (N759)? data_n_45__8_ : 
                      (N761)? data_n_46__8_ : 
                      (N763)? data_n_47__8_ : 
                      (N765)? data_n_48__8_ : 
                      (N767)? data_n_49__8_ : 
                      (N769)? data_n_50__8_ : 
                      (N771)? data_n_51__8_ : 
                      (N773)? data_n_52__8_ : 
                      (N775)? data_n_53__8_ : 
                      (N777)? data_n_54__8_ : 
                      (N779)? data_n_55__8_ : 
                      (N781)? data_n_56__8_ : 
                      (N783)? data_n_57__8_ : 
                      (N785)? data_n_58__8_ : 
                      (N787)? data_n_59__8_ : 
                      (N789)? data_n_60__8_ : 
                      (N791)? data_n_61__8_ : 
                      (N793)? data_n_62__8_ : 
                      (N795)? data_n_63__8_ : 1'b0;
  assign data_nn[7] = (N732)? data_o[7] : 
                      (N734)? data_o[23] : 
                      (N736)? data_o[39] : 
                      (N738)? data_o[55] : 
                      (N740)? data_o[71] : 
                      (N742)? data_o[87] : 
                      (N744)? data_o[103] : 
                      (N746)? data_o[119] : 
                      (N748)? data_o[135] : 
                      (N750)? data_o[151] : 
                      (N752)? data_o[167] : 
                      (N754)? data_o[183] : 
                      (N756)? data_o[199] : 
                      (N758)? data_o[215] : 
                      (N760)? data_o[231] : 
                      (N762)? data_o[247] : 
                      (N764)? data_o[263] : 
                      (N766)? data_o[279] : 
                      (N768)? data_o[295] : 
                      (N770)? data_o[311] : 
                      (N772)? data_o[327] : 
                      (N774)? data_o[343] : 
                      (N776)? data_o[359] : 
                      (N778)? data_o[375] : 
                      (N780)? data_o[391] : 
                      (N782)? data_o[407] : 
                      (N784)? data_o[423] : 
                      (N786)? data_o[439] : 
                      (N788)? data_o[455] : 
                      (N790)? data_o[471] : 
                      (N792)? data_o[487] : 
                      (N794)? data_o[503] : 
                      (N733)? data_n_32__7_ : 
                      (N735)? data_n_33__7_ : 
                      (N737)? data_n_34__7_ : 
                      (N739)? data_n_35__7_ : 
                      (N741)? data_n_36__7_ : 
                      (N743)? data_n_37__7_ : 
                      (N745)? data_n_38__7_ : 
                      (N747)? data_n_39__7_ : 
                      (N749)? data_n_40__7_ : 
                      (N751)? data_n_41__7_ : 
                      (N753)? data_n_42__7_ : 
                      (N755)? data_n_43__7_ : 
                      (N757)? data_n_44__7_ : 
                      (N759)? data_n_45__7_ : 
                      (N761)? data_n_46__7_ : 
                      (N763)? data_n_47__7_ : 
                      (N765)? data_n_48__7_ : 
                      (N767)? data_n_49__7_ : 
                      (N769)? data_n_50__7_ : 
                      (N771)? data_n_51__7_ : 
                      (N773)? data_n_52__7_ : 
                      (N775)? data_n_53__7_ : 
                      (N777)? data_n_54__7_ : 
                      (N779)? data_n_55__7_ : 
                      (N781)? data_n_56__7_ : 
                      (N783)? data_n_57__7_ : 
                      (N785)? data_n_58__7_ : 
                      (N787)? data_n_59__7_ : 
                      (N789)? data_n_60__7_ : 
                      (N791)? data_n_61__7_ : 
                      (N793)? data_n_62__7_ : 
                      (N795)? data_n_63__7_ : 1'b0;
  assign data_nn[6] = (N732)? data_o[6] : 
                      (N734)? data_o[22] : 
                      (N736)? data_o[38] : 
                      (N738)? data_o[54] : 
                      (N740)? data_o[70] : 
                      (N742)? data_o[86] : 
                      (N744)? data_o[102] : 
                      (N746)? data_o[118] : 
                      (N748)? data_o[134] : 
                      (N750)? data_o[150] : 
                      (N752)? data_o[166] : 
                      (N754)? data_o[182] : 
                      (N756)? data_o[198] : 
                      (N758)? data_o[214] : 
                      (N760)? data_o[230] : 
                      (N762)? data_o[246] : 
                      (N764)? data_o[262] : 
                      (N766)? data_o[278] : 
                      (N768)? data_o[294] : 
                      (N770)? data_o[310] : 
                      (N772)? data_o[326] : 
                      (N774)? data_o[342] : 
                      (N776)? data_o[358] : 
                      (N778)? data_o[374] : 
                      (N780)? data_o[390] : 
                      (N782)? data_o[406] : 
                      (N784)? data_o[422] : 
                      (N786)? data_o[438] : 
                      (N788)? data_o[454] : 
                      (N790)? data_o[470] : 
                      (N792)? data_o[486] : 
                      (N794)? data_o[502] : 
                      (N733)? data_n_32__6_ : 
                      (N735)? data_n_33__6_ : 
                      (N737)? data_n_34__6_ : 
                      (N739)? data_n_35__6_ : 
                      (N741)? data_n_36__6_ : 
                      (N743)? data_n_37__6_ : 
                      (N745)? data_n_38__6_ : 
                      (N747)? data_n_39__6_ : 
                      (N749)? data_n_40__6_ : 
                      (N751)? data_n_41__6_ : 
                      (N753)? data_n_42__6_ : 
                      (N755)? data_n_43__6_ : 
                      (N757)? data_n_44__6_ : 
                      (N759)? data_n_45__6_ : 
                      (N761)? data_n_46__6_ : 
                      (N763)? data_n_47__6_ : 
                      (N765)? data_n_48__6_ : 
                      (N767)? data_n_49__6_ : 
                      (N769)? data_n_50__6_ : 
                      (N771)? data_n_51__6_ : 
                      (N773)? data_n_52__6_ : 
                      (N775)? data_n_53__6_ : 
                      (N777)? data_n_54__6_ : 
                      (N779)? data_n_55__6_ : 
                      (N781)? data_n_56__6_ : 
                      (N783)? data_n_57__6_ : 
                      (N785)? data_n_58__6_ : 
                      (N787)? data_n_59__6_ : 
                      (N789)? data_n_60__6_ : 
                      (N791)? data_n_61__6_ : 
                      (N793)? data_n_62__6_ : 
                      (N795)? data_n_63__6_ : 1'b0;
  assign data_nn[5] = (N732)? data_o[5] : 
                      (N734)? data_o[21] : 
                      (N736)? data_o[37] : 
                      (N738)? data_o[53] : 
                      (N740)? data_o[69] : 
                      (N742)? data_o[85] : 
                      (N744)? data_o[101] : 
                      (N746)? data_o[117] : 
                      (N748)? data_o[133] : 
                      (N750)? data_o[149] : 
                      (N752)? data_o[165] : 
                      (N754)? data_o[181] : 
                      (N756)? data_o[197] : 
                      (N758)? data_o[213] : 
                      (N760)? data_o[229] : 
                      (N762)? data_o[245] : 
                      (N764)? data_o[261] : 
                      (N766)? data_o[277] : 
                      (N768)? data_o[293] : 
                      (N770)? data_o[309] : 
                      (N772)? data_o[325] : 
                      (N774)? data_o[341] : 
                      (N776)? data_o[357] : 
                      (N778)? data_o[373] : 
                      (N780)? data_o[389] : 
                      (N782)? data_o[405] : 
                      (N784)? data_o[421] : 
                      (N786)? data_o[437] : 
                      (N788)? data_o[453] : 
                      (N790)? data_o[469] : 
                      (N792)? data_o[485] : 
                      (N794)? data_o[501] : 
                      (N733)? data_n_32__5_ : 
                      (N735)? data_n_33__5_ : 
                      (N737)? data_n_34__5_ : 
                      (N739)? data_n_35__5_ : 
                      (N741)? data_n_36__5_ : 
                      (N743)? data_n_37__5_ : 
                      (N745)? data_n_38__5_ : 
                      (N747)? data_n_39__5_ : 
                      (N749)? data_n_40__5_ : 
                      (N751)? data_n_41__5_ : 
                      (N753)? data_n_42__5_ : 
                      (N755)? data_n_43__5_ : 
                      (N757)? data_n_44__5_ : 
                      (N759)? data_n_45__5_ : 
                      (N761)? data_n_46__5_ : 
                      (N763)? data_n_47__5_ : 
                      (N765)? data_n_48__5_ : 
                      (N767)? data_n_49__5_ : 
                      (N769)? data_n_50__5_ : 
                      (N771)? data_n_51__5_ : 
                      (N773)? data_n_52__5_ : 
                      (N775)? data_n_53__5_ : 
                      (N777)? data_n_54__5_ : 
                      (N779)? data_n_55__5_ : 
                      (N781)? data_n_56__5_ : 
                      (N783)? data_n_57__5_ : 
                      (N785)? data_n_58__5_ : 
                      (N787)? data_n_59__5_ : 
                      (N789)? data_n_60__5_ : 
                      (N791)? data_n_61__5_ : 
                      (N793)? data_n_62__5_ : 
                      (N795)? data_n_63__5_ : 1'b0;
  assign data_nn[4] = (N732)? data_o[4] : 
                      (N734)? data_o[20] : 
                      (N736)? data_o[36] : 
                      (N738)? data_o[52] : 
                      (N740)? data_o[68] : 
                      (N742)? data_o[84] : 
                      (N744)? data_o[100] : 
                      (N746)? data_o[116] : 
                      (N748)? data_o[132] : 
                      (N750)? data_o[148] : 
                      (N752)? data_o[164] : 
                      (N754)? data_o[180] : 
                      (N756)? data_o[196] : 
                      (N758)? data_o[212] : 
                      (N760)? data_o[228] : 
                      (N762)? data_o[244] : 
                      (N764)? data_o[260] : 
                      (N766)? data_o[276] : 
                      (N768)? data_o[292] : 
                      (N770)? data_o[308] : 
                      (N772)? data_o[324] : 
                      (N774)? data_o[340] : 
                      (N776)? data_o[356] : 
                      (N778)? data_o[372] : 
                      (N780)? data_o[388] : 
                      (N782)? data_o[404] : 
                      (N784)? data_o[420] : 
                      (N786)? data_o[436] : 
                      (N788)? data_o[452] : 
                      (N790)? data_o[468] : 
                      (N792)? data_o[484] : 
                      (N794)? data_o[500] : 
                      (N733)? data_n_32__4_ : 
                      (N735)? data_n_33__4_ : 
                      (N737)? data_n_34__4_ : 
                      (N739)? data_n_35__4_ : 
                      (N741)? data_n_36__4_ : 
                      (N743)? data_n_37__4_ : 
                      (N745)? data_n_38__4_ : 
                      (N747)? data_n_39__4_ : 
                      (N749)? data_n_40__4_ : 
                      (N751)? data_n_41__4_ : 
                      (N753)? data_n_42__4_ : 
                      (N755)? data_n_43__4_ : 
                      (N757)? data_n_44__4_ : 
                      (N759)? data_n_45__4_ : 
                      (N761)? data_n_46__4_ : 
                      (N763)? data_n_47__4_ : 
                      (N765)? data_n_48__4_ : 
                      (N767)? data_n_49__4_ : 
                      (N769)? data_n_50__4_ : 
                      (N771)? data_n_51__4_ : 
                      (N773)? data_n_52__4_ : 
                      (N775)? data_n_53__4_ : 
                      (N777)? data_n_54__4_ : 
                      (N779)? data_n_55__4_ : 
                      (N781)? data_n_56__4_ : 
                      (N783)? data_n_57__4_ : 
                      (N785)? data_n_58__4_ : 
                      (N787)? data_n_59__4_ : 
                      (N789)? data_n_60__4_ : 
                      (N791)? data_n_61__4_ : 
                      (N793)? data_n_62__4_ : 
                      (N795)? data_n_63__4_ : 1'b0;
  assign data_nn[3] = (N732)? data_o[3] : 
                      (N734)? data_o[19] : 
                      (N736)? data_o[35] : 
                      (N738)? data_o[51] : 
                      (N740)? data_o[67] : 
                      (N742)? data_o[83] : 
                      (N744)? data_o[99] : 
                      (N746)? data_o[115] : 
                      (N748)? data_o[131] : 
                      (N750)? data_o[147] : 
                      (N752)? data_o[163] : 
                      (N754)? data_o[179] : 
                      (N756)? data_o[195] : 
                      (N758)? data_o[211] : 
                      (N760)? data_o[227] : 
                      (N762)? data_o[243] : 
                      (N764)? data_o[259] : 
                      (N766)? data_o[275] : 
                      (N768)? data_o[291] : 
                      (N770)? data_o[307] : 
                      (N772)? data_o[323] : 
                      (N774)? data_o[339] : 
                      (N776)? data_o[355] : 
                      (N778)? data_o[371] : 
                      (N780)? data_o[387] : 
                      (N782)? data_o[403] : 
                      (N784)? data_o[419] : 
                      (N786)? data_o[435] : 
                      (N788)? data_o[451] : 
                      (N790)? data_o[467] : 
                      (N792)? data_o[483] : 
                      (N794)? data_o[499] : 
                      (N733)? data_n_32__3_ : 
                      (N735)? data_n_33__3_ : 
                      (N737)? data_n_34__3_ : 
                      (N739)? data_n_35__3_ : 
                      (N741)? data_n_36__3_ : 
                      (N743)? data_n_37__3_ : 
                      (N745)? data_n_38__3_ : 
                      (N747)? data_n_39__3_ : 
                      (N749)? data_n_40__3_ : 
                      (N751)? data_n_41__3_ : 
                      (N753)? data_n_42__3_ : 
                      (N755)? data_n_43__3_ : 
                      (N757)? data_n_44__3_ : 
                      (N759)? data_n_45__3_ : 
                      (N761)? data_n_46__3_ : 
                      (N763)? data_n_47__3_ : 
                      (N765)? data_n_48__3_ : 
                      (N767)? data_n_49__3_ : 
                      (N769)? data_n_50__3_ : 
                      (N771)? data_n_51__3_ : 
                      (N773)? data_n_52__3_ : 
                      (N775)? data_n_53__3_ : 
                      (N777)? data_n_54__3_ : 
                      (N779)? data_n_55__3_ : 
                      (N781)? data_n_56__3_ : 
                      (N783)? data_n_57__3_ : 
                      (N785)? data_n_58__3_ : 
                      (N787)? data_n_59__3_ : 
                      (N789)? data_n_60__3_ : 
                      (N791)? data_n_61__3_ : 
                      (N793)? data_n_62__3_ : 
                      (N795)? data_n_63__3_ : 1'b0;
  assign data_nn[2] = (N732)? data_o[2] : 
                      (N734)? data_o[18] : 
                      (N736)? data_o[34] : 
                      (N738)? data_o[50] : 
                      (N740)? data_o[66] : 
                      (N742)? data_o[82] : 
                      (N744)? data_o[98] : 
                      (N746)? data_o[114] : 
                      (N748)? data_o[130] : 
                      (N750)? data_o[146] : 
                      (N752)? data_o[162] : 
                      (N754)? data_o[178] : 
                      (N756)? data_o[194] : 
                      (N758)? data_o[210] : 
                      (N760)? data_o[226] : 
                      (N762)? data_o[242] : 
                      (N764)? data_o[258] : 
                      (N766)? data_o[274] : 
                      (N768)? data_o[290] : 
                      (N770)? data_o[306] : 
                      (N772)? data_o[322] : 
                      (N774)? data_o[338] : 
                      (N776)? data_o[354] : 
                      (N778)? data_o[370] : 
                      (N780)? data_o[386] : 
                      (N782)? data_o[402] : 
                      (N784)? data_o[418] : 
                      (N786)? data_o[434] : 
                      (N788)? data_o[450] : 
                      (N790)? data_o[466] : 
                      (N792)? data_o[482] : 
                      (N794)? data_o[498] : 
                      (N733)? data_n_32__2_ : 
                      (N735)? data_n_33__2_ : 
                      (N737)? data_n_34__2_ : 
                      (N739)? data_n_35__2_ : 
                      (N741)? data_n_36__2_ : 
                      (N743)? data_n_37__2_ : 
                      (N745)? data_n_38__2_ : 
                      (N747)? data_n_39__2_ : 
                      (N749)? data_n_40__2_ : 
                      (N751)? data_n_41__2_ : 
                      (N753)? data_n_42__2_ : 
                      (N755)? data_n_43__2_ : 
                      (N757)? data_n_44__2_ : 
                      (N759)? data_n_45__2_ : 
                      (N761)? data_n_46__2_ : 
                      (N763)? data_n_47__2_ : 
                      (N765)? data_n_48__2_ : 
                      (N767)? data_n_49__2_ : 
                      (N769)? data_n_50__2_ : 
                      (N771)? data_n_51__2_ : 
                      (N773)? data_n_52__2_ : 
                      (N775)? data_n_53__2_ : 
                      (N777)? data_n_54__2_ : 
                      (N779)? data_n_55__2_ : 
                      (N781)? data_n_56__2_ : 
                      (N783)? data_n_57__2_ : 
                      (N785)? data_n_58__2_ : 
                      (N787)? data_n_59__2_ : 
                      (N789)? data_n_60__2_ : 
                      (N791)? data_n_61__2_ : 
                      (N793)? data_n_62__2_ : 
                      (N795)? data_n_63__2_ : 1'b0;
  assign data_nn[1] = (N732)? data_o[1] : 
                      (N734)? data_o[17] : 
                      (N736)? data_o[33] : 
                      (N738)? data_o[49] : 
                      (N740)? data_o[65] : 
                      (N742)? data_o[81] : 
                      (N744)? data_o[97] : 
                      (N746)? data_o[113] : 
                      (N748)? data_o[129] : 
                      (N750)? data_o[145] : 
                      (N752)? data_o[161] : 
                      (N754)? data_o[177] : 
                      (N756)? data_o[193] : 
                      (N758)? data_o[209] : 
                      (N760)? data_o[225] : 
                      (N762)? data_o[241] : 
                      (N764)? data_o[257] : 
                      (N766)? data_o[273] : 
                      (N768)? data_o[289] : 
                      (N770)? data_o[305] : 
                      (N772)? data_o[321] : 
                      (N774)? data_o[337] : 
                      (N776)? data_o[353] : 
                      (N778)? data_o[369] : 
                      (N780)? data_o[385] : 
                      (N782)? data_o[401] : 
                      (N784)? data_o[417] : 
                      (N786)? data_o[433] : 
                      (N788)? data_o[449] : 
                      (N790)? data_o[465] : 
                      (N792)? data_o[481] : 
                      (N794)? data_o[497] : 
                      (N733)? data_n_32__1_ : 
                      (N735)? data_n_33__1_ : 
                      (N737)? data_n_34__1_ : 
                      (N739)? data_n_35__1_ : 
                      (N741)? data_n_36__1_ : 
                      (N743)? data_n_37__1_ : 
                      (N745)? data_n_38__1_ : 
                      (N747)? data_n_39__1_ : 
                      (N749)? data_n_40__1_ : 
                      (N751)? data_n_41__1_ : 
                      (N753)? data_n_42__1_ : 
                      (N755)? data_n_43__1_ : 
                      (N757)? data_n_44__1_ : 
                      (N759)? data_n_45__1_ : 
                      (N761)? data_n_46__1_ : 
                      (N763)? data_n_47__1_ : 
                      (N765)? data_n_48__1_ : 
                      (N767)? data_n_49__1_ : 
                      (N769)? data_n_50__1_ : 
                      (N771)? data_n_51__1_ : 
                      (N773)? data_n_52__1_ : 
                      (N775)? data_n_53__1_ : 
                      (N777)? data_n_54__1_ : 
                      (N779)? data_n_55__1_ : 
                      (N781)? data_n_56__1_ : 
                      (N783)? data_n_57__1_ : 
                      (N785)? data_n_58__1_ : 
                      (N787)? data_n_59__1_ : 
                      (N789)? data_n_60__1_ : 
                      (N791)? data_n_61__1_ : 
                      (N793)? data_n_62__1_ : 
                      (N795)? data_n_63__1_ : 1'b0;
  assign data_nn[0] = (N732)? data_o[0] : 
                      (N734)? data_o[16] : 
                      (N736)? data_o[32] : 
                      (N738)? data_o[48] : 
                      (N740)? data_o[64] : 
                      (N742)? data_o[80] : 
                      (N744)? data_o[96] : 
                      (N746)? data_o[112] : 
                      (N748)? data_o[128] : 
                      (N750)? data_o[144] : 
                      (N752)? data_o[160] : 
                      (N754)? data_o[176] : 
                      (N756)? data_o[192] : 
                      (N758)? data_o[208] : 
                      (N760)? data_o[224] : 
                      (N762)? data_o[240] : 
                      (N764)? data_o[256] : 
                      (N766)? data_o[272] : 
                      (N768)? data_o[288] : 
                      (N770)? data_o[304] : 
                      (N772)? data_o[320] : 
                      (N774)? data_o[336] : 
                      (N776)? data_o[352] : 
                      (N778)? data_o[368] : 
                      (N780)? data_o[384] : 
                      (N782)? data_o[400] : 
                      (N784)? data_o[416] : 
                      (N786)? data_o[432] : 
                      (N788)? data_o[448] : 
                      (N790)? data_o[464] : 
                      (N792)? data_o[480] : 
                      (N794)? data_o[496] : 
                      (N733)? data_n_32__0_ : 
                      (N735)? data_n_33__0_ : 
                      (N737)? data_n_34__0_ : 
                      (N739)? data_n_35__0_ : 
                      (N741)? data_n_36__0_ : 
                      (N743)? data_n_37__0_ : 
                      (N745)? data_n_38__0_ : 
                      (N747)? data_n_39__0_ : 
                      (N749)? data_n_40__0_ : 
                      (N751)? data_n_41__0_ : 
                      (N753)? data_n_42__0_ : 
                      (N755)? data_n_43__0_ : 
                      (N757)? data_n_44__0_ : 
                      (N759)? data_n_45__0_ : 
                      (N761)? data_n_46__0_ : 
                      (N763)? data_n_47__0_ : 
                      (N765)? data_n_48__0_ : 
                      (N767)? data_n_49__0_ : 
                      (N769)? data_n_50__0_ : 
                      (N771)? data_n_51__0_ : 
                      (N773)? data_n_52__0_ : 
                      (N775)? data_n_53__0_ : 
                      (N777)? data_n_54__0_ : 
                      (N779)? data_n_55__0_ : 
                      (N781)? data_n_56__0_ : 
                      (N783)? data_n_57__0_ : 
                      (N785)? data_n_58__0_ : 
                      (N787)? data_n_59__0_ : 
                      (N789)? data_n_60__0_ : 
                      (N791)? data_n_61__0_ : 
                      (N793)? data_n_62__0_ : 
                      (N795)? data_n_63__0_ : 1'b0;
  assign { N408, N407, N406, N405, N404, N403 } = num_els_r + N402;
  assign num_els_n = { N408, N407, N406, N405, N404, N403 } - yumi_cnt_i;
  assign N1205 = ~num_els_r[5];
  assign N1206 = num_els_r[3] & num_els_r[4];
  assign N1207 = N0 & num_els_r[4];
  assign N0 = ~num_els_r[3];
  assign N1208 = num_els_r[3] & N1;
  assign N1 = ~num_els_r[4];
  assign N1209 = N2 & N3;
  assign N2 = ~num_els_r[3];
  assign N3 = ~num_els_r[4];
  assign N1210 = num_els_r[5] & N1206;
  assign N1211 = num_els_r[5] & N1207;
  assign N1212 = num_els_r[5] & N1208;
  assign N1213 = num_els_r[5] & N1209;
  assign N1214 = N1205 & N1206;
  assign N1215 = N1205 & N1207;
  assign N1216 = N1205 & N1208;
  assign N1217 = N1205 & N1209;
  assign N1218 = ~num_els_r[2];
  assign N1219 = num_els_r[0] & num_els_r[1];
  assign N1220 = N4 & num_els_r[1];
  assign N4 = ~num_els_r[0];
  assign N1221 = num_els_r[0] & N5;
  assign N5 = ~num_els_r[1];
  assign N1222 = N6 & N7;
  assign N6 = ~num_els_r[0];
  assign N7 = ~num_els_r[1];
  assign N1223 = num_els_r[2] & N1219;
  assign N1224 = num_els_r[2] & N1220;
  assign N1225 = num_els_r[2] & N1221;
  assign N1226 = num_els_r[2] & N1222;
  assign N1227 = N1218 & N1219;
  assign N1228 = N1218 & N1220;
  assign N1229 = N1218 & N1221;
  assign N1230 = N1218 & N1222;
  assign N472 = N1210 & N1223;
  assign N471 = N1210 & N1224;
  assign N470 = N1210 & N1225;
  assign N469 = N1210 & N1226;
  assign N468 = N1210 & N1227;
  assign N467 = N1210 & N1228;
  assign N466 = N1210 & N1229;
  assign N465 = N1210 & N1230;
  assign N464 = N1211 & N1223;
  assign N463 = N1211 & N1224;
  assign N462 = N1211 & N1225;
  assign N461 = N1211 & N1226;
  assign N460 = N1211 & N1227;
  assign N459 = N1211 & N1228;
  assign N458 = N1211 & N1229;
  assign N457 = N1211 & N1230;
  assign N456 = N1212 & N1223;
  assign N455 = N1212 & N1224;
  assign N454 = N1212 & N1225;
  assign N453 = N1212 & N1226;
  assign N452 = N1212 & N1227;
  assign N451 = N1212 & N1228;
  assign N450 = N1212 & N1229;
  assign N449 = N1212 & N1230;
  assign N448 = N1213 & N1223;
  assign N447 = N1213 & N1224;
  assign N446 = N1213 & N1225;
  assign N445 = N1213 & N1226;
  assign N444 = N1213 & N1227;
  assign N443 = N1213 & N1228;
  assign N442 = N1213 & N1229;
  assign N441 = N1213 & N1230;
  assign N440 = N1214 & N1223;
  assign N439 = N1214 & N1224;
  assign N438 = N1214 & N1225;
  assign N437 = N1214 & N1226;
  assign N436 = N1214 & N1227;
  assign N435 = N1214 & N1228;
  assign N434 = N1214 & N1229;
  assign N433 = N1214 & N1230;
  assign N432 = N1215 & N1223;
  assign N431 = N1215 & N1224;
  assign N430 = N1215 & N1225;
  assign N429 = N1215 & N1226;
  assign N428 = N1215 & N1227;
  assign N427 = N1215 & N1228;
  assign N426 = N1215 & N1229;
  assign N425 = N1215 & N1230;
  assign N424 = N1216 & N1223;
  assign N423 = N1216 & N1224;
  assign N422 = N1216 & N1225;
  assign N421 = N1216 & N1226;
  assign N420 = N1216 & N1227;
  assign N419 = N1216 & N1228;
  assign N418 = N1216 & N1229;
  assign N417 = N1216 & N1230;
  assign N416 = N1217 & N1223;
  assign N415 = N1217 & N1224;
  assign N414 = N1217 & N1225;
  assign N413 = N1217 & N1226;
  assign N412 = N1217 & N1227;
  assign N411 = N1217 & N1228;
  assign N410 = N1217 & N1229;
  assign N409 = N1217 & N1230;
  assign N1231 = num_els_r[3] & num_els_r[4];
  assign N1232 = N8 & num_els_r[4];
  assign N8 = ~num_els_r[3];
  assign N1233 = num_els_r[3] & N9;
  assign N9 = ~num_els_r[4];
  assign N1234 = N10 & N11;
  assign N10 = ~num_els_r[3];
  assign N11 = ~num_els_r[4];
  assign N1235 = num_els_r[5] & N1231;
  assign N1236 = num_els_r[5] & N1232;
  assign N1237 = num_els_r[5] & N1233;
  assign N1238 = num_els_r[5] & N1234;
  assign N1239 = N1205 & N1231;
  assign N1240 = N1205 & N1232;
  assign N1241 = N1205 & N1233;
  assign N1242 = N1205 & N1234;
  assign N1243 = num_els_r[0] & num_els_r[1];
  assign N1244 = N12 & num_els_r[1];
  assign N12 = ~num_els_r[0];
  assign N1245 = num_els_r[0] & N13;
  assign N13 = ~num_els_r[1];
  assign N1246 = N14 & N15;
  assign N14 = ~num_els_r[0];
  assign N15 = ~num_els_r[1];
  assign N1247 = num_els_r[2] & N1243;
  assign N1248 = num_els_r[2] & N1244;
  assign N1249 = num_els_r[2] & N1245;
  assign N1250 = num_els_r[2] & N1246;
  assign N1251 = N1218 & N1243;
  assign N1252 = N1218 & N1244;
  assign N1253 = N1218 & N1245;
  assign N1254 = N1218 & N1246;
  assign N600 = N1235 & N1247;
  assign N599 = N1235 & N1248;
  assign N598 = N1235 & N1249;
  assign N597 = N1235 & N1250;
  assign N596 = N1235 & N1251;
  assign N595 = N1235 & N1252;
  assign N594 = N1235 & N1253;
  assign N593 = N1235 & N1254;
  assign N592 = N1236 & N1247;
  assign N591 = N1236 & N1248;
  assign N590 = N1236 & N1249;
  assign N589 = N1236 & N1250;
  assign N588 = N1236 & N1251;
  assign N587 = N1236 & N1252;
  assign N586 = N1236 & N1253;
  assign N585 = N1236 & N1254;
  assign N584 = N1237 & N1247;
  assign N583 = N1237 & N1248;
  assign N582 = N1237 & N1249;
  assign N581 = N1237 & N1250;
  assign N580 = N1237 & N1251;
  assign N579 = N1237 & N1252;
  assign N578 = N1237 & N1253;
  assign N577 = N1237 & N1254;
  assign N576 = N1238 & N1247;
  assign N575 = N1238 & N1248;
  assign N574 = N1238 & N1249;
  assign N573 = N1238 & N1250;
  assign N572 = N1238 & N1251;
  assign N571 = N1238 & N1252;
  assign N570 = N1238 & N1253;
  assign N569 = N1238 & N1254;
  assign N568 = N1239 & N1247;
  assign N567 = N1239 & N1248;
  assign N566 = N1239 & N1249;
  assign N565 = N1239 & N1250;
  assign N564 = N1239 & N1251;
  assign N563 = N1239 & N1252;
  assign N562 = N1239 & N1253;
  assign N561 = N1239 & N1254;
  assign N560 = N1240 & N1247;
  assign N559 = N1240 & N1248;
  assign N558 = N1240 & N1249;
  assign N557 = N1240 & N1250;
  assign N556 = N1240 & N1251;
  assign N555 = N1240 & N1252;
  assign N554 = N1240 & N1253;
  assign N553 = N1240 & N1254;
  assign N552 = N1241 & N1247;
  assign N551 = N1241 & N1248;
  assign N550 = N1241 & N1249;
  assign N549 = N1241 & N1250;
  assign N548 = N1241 & N1251;
  assign N547 = N1241 & N1252;
  assign N546 = N1241 & N1253;
  assign N545 = N1241 & N1254;
  assign N544 = N1242 & N1247;
  assign N543 = N1242 & N1248;
  assign N542 = N1242 & N1249;
  assign N541 = N1242 & N1250;
  assign N540 = N1242 & N1251;
  assign N539 = N1242 & N1252;
  assign N538 = N1242 & N1253;
  assign N537 = N1242 & N1254;
  assign N1255 = ~yumi_cnt_i[5];
  assign N1256 = N1255 & N1319;
  assign N1257 = N1255 & N1320;
  assign N1258 = N1255 & N1321;
  assign N1259 = N1255 & N1322;
  assign N1260 = ~yumi_cnt_i[2];
  assign N1261 = N1260 & N1331;
  assign N1262 = N1260 & N1332;
  assign N1263 = N1260 & N1333;
  assign N1264 = N1260 & N1334;
  assign N1265 = N1323 & N1261;
  assign N1266 = N1323 & N1262;
  assign N841 = N1323 & N1263;
  assign N840 = N1323 & N1264;
  assign N839 = N1324 & N1261;
  assign N838 = N1324 & N1262;
  assign N837 = N1324 & N1263;
  assign N836 = N1324 & N1264;
  assign N835 = N1325 & N1261;
  assign N834 = N1325 & N1262;
  assign N833 = N1325 & N1263;
  assign N832 = N1325 & N1264;
  assign N831 = N1326 & N1261;
  assign N830 = N1326 & N1262;
  assign N829 = N1326 & N1263;
  assign N828 = N1326 & N1264;
  assign N827 = N1256 & N1335;
  assign N826 = N1256 & N1336;
  assign N825 = N1256 & N1337;
  assign N824 = N1256 & N1338;
  assign N823 = N1256 & N1261;
  assign N822 = N1256 & N1262;
  assign N821 = N1256 & N1263;
  assign N820 = N1256 & N1264;
  assign N819 = N1257 & N1335;
  assign N818 = N1257 & N1336;
  assign N817 = N1257 & N1337;
  assign N816 = N1257 & N1338;
  assign N815 = N1257 & N1261;
  assign N814 = N1257 & N1262;
  assign N813 = N1257 & N1263;
  assign N812 = N1257 & N1264;
  assign N811 = N1258 & N1335;
  assign N810 = N1258 & N1336;
  assign N809 = N1258 & N1337;
  assign N808 = N1258 & N1338;
  assign N807 = N1258 & N1261;
  assign N806 = N1258 & N1262;
  assign N805 = N1258 & N1263;
  assign N804 = N1258 & N1264;
  assign N803 = N1259 & N1335;
  assign N802 = N1259 & N1336;
  assign N801 = N1259 & N1337;
  assign N800 = N1259 & N1338;
  assign N799 = N1259 & N1261;
  assign N798 = N1259 & N1262;
  assign N797 = N1259 & N1263;
  assign N796 = N1259 & N1264;
  assign N1267 = N1290 & N1339;
  assign N1268 = N1290 & N1340;
  assign N1269 = N1290 & N1341;
  assign N1270 = N1290 & N1342;
  assign N865 = N1291 & N1339;
  assign N864 = N1291 & N1340;
  assign N863 = N1291 & N1341;
  assign N862 = N1291 & N1342;
  assign N861 = N1292 & N1339;
  assign N860 = N1292 & N1340;
  assign N859 = N1292 & N1341;
  assign N858 = N1292 & N1342;
  assign N857 = N1327 & N1297;
  assign N856 = N1327 & N1298;
  assign N855 = N1327 & N1299;
  assign N854 = N1327 & N1300;
  assign N853 = N1328 & N1297;
  assign N852 = N1328 & N1298;
  assign N851 = N1328 & N1299;
  assign N850 = N1328 & N1300;
  assign N849 = N1329 & N1297;
  assign N848 = N1329 & N1298;
  assign N847 = N1329 & N1299;
  assign N846 = N1329 & N1300;
  assign N845 = N1330 & N1297;
  assign N844 = N1330 & N1298;
  assign N843 = N1330 & N1299;
  assign N842 = N1330 & N1300;
  assign N1271 = N1272 & N1304;
  assign N885 = N1273 & N1301;
  assign N884 = N1273 & N1302;
  assign N883 = N1273 & N1303;
  assign N882 = N1273 & N1304;
  assign N881 = N1293 & N1278;
  assign N880 = N1293 & N1279;
  assign N879 = N1293 & N1280;
  assign N878 = N1293 & N1281;
  assign N877 = N1294 & N1278;
  assign N876 = N1294 & N1279;
  assign N875 = N1294 & N1280;
  assign N874 = N1294 & N1281;
  assign N873 = N1295 & N1278;
  assign N872 = N1295 & N1279;
  assign N871 = N1295 & N1280;
  assign N870 = N1295 & N1281;
  assign N869 = N1296 & N1278;
  assign N868 = N1296 & N1279;
  assign N867 = N1296 & N1280;
  assign N866 = N1296 & N1281;
  assign N1272 = yumi_cnt_i[5] & N1321;
  assign N1273 = yumi_cnt_i[5] & N1322;
  assign N1274 = N1255 & N1319;
  assign N1275 = N1255 & N1320;
  assign N1276 = N1255 & N1321;
  assign N1277 = N1255 & N1322;
  assign N1278 = yumi_cnt_i[2] & N1331;
  assign N1279 = yumi_cnt_i[2] & N1332;
  assign N1280 = yumi_cnt_i[2] & N1333;
  assign N1281 = yumi_cnt_i[2] & N1334;
  assign N1282 = N1260 & N1331;
  assign N1283 = N1260 & N1332;
  assign N1284 = N1260 & N1333;
  assign N1285 = N1260 & N1334;
  assign N1286 = N1273 & N1278;
  assign N1287 = N1273 & N1279;
  assign N1288 = N1273 & N1280;
  assign N1289 = N1273 & N1281;
  assign N920 = N1273 & N1283;
  assign N919 = N1273 & N1284;
  assign N918 = N1273 & N1285;
  assign N917 = N1274 & N1278;
  assign N916 = N1274 & N1279;
  assign N915 = N1274 & N1280;
  assign N914 = N1274 & N1281;
  assign N913 = N1274 & N1282;
  assign N912 = N1274 & N1283;
  assign N911 = N1274 & N1284;
  assign N910 = N1274 & N1285;
  assign N909 = N1275 & N1278;
  assign N908 = N1275 & N1279;
  assign N907 = N1275 & N1280;
  assign N906 = N1275 & N1281;
  assign N905 = N1275 & N1282;
  assign N904 = N1275 & N1283;
  assign N903 = N1275 & N1284;
  assign N902 = N1275 & N1285;
  assign N901 = N1276 & N1278;
  assign N900 = N1276 & N1279;
  assign N899 = N1276 & N1280;
  assign N898 = N1276 & N1281;
  assign N897 = N1276 & N1282;
  assign N896 = N1276 & N1283;
  assign N895 = N1276 & N1284;
  assign N894 = N1276 & N1285;
  assign N893 = N1277 & N1278;
  assign N892 = N1277 & N1279;
  assign N891 = N1277 & N1280;
  assign N890 = N1277 & N1281;
  assign N889 = N1277 & N1282;
  assign N888 = N1277 & N1283;
  assign N887 = N1277 & N1284;
  assign N886 = N1277 & N1285;
  assign N1290 = yumi_cnt_i[5] & N1320;
  assign N1291 = yumi_cnt_i[5] & N1321;
  assign N1292 = yumi_cnt_i[5] & N1322;
  assign N1293 = N1255 & N1319;
  assign N1294 = N1255 & N1320;
  assign N1295 = N1255 & N1321;
  assign N1296 = N1255 & N1322;
  assign N1297 = yumi_cnt_i[2] & N1331;
  assign N1298 = yumi_cnt_i[2] & N1332;
  assign N1299 = yumi_cnt_i[2] & N1333;
  assign N1300 = yumi_cnt_i[2] & N1334;
  assign N1301 = N1260 & N1331;
  assign N1302 = N1260 & N1332;
  assign N1303 = N1260 & N1333;
  assign N1304 = N1260 & N1334;
  assign N1305 = N1291 & N1297;
  assign N1306 = N1291 & N1298;
  assign N1307 = N1291 & N1299;
  assign N1308 = N1291 & N1300;
  assign N1309 = N1291 & N1301;
  assign N1310 = N1291 & N1302;
  assign N1311 = N1291 & N1303;
  assign N1312 = N1291 & N1304;
  assign N1313 = N1292 & N1297;
  assign N1314 = N1292 & N1298;
  assign N1315 = N1292 & N1299;
  assign N1316 = N1292 & N1300;
  assign N1317 = N1292 & N1301;
  assign N1318 = N1292 & N1302;
  assign N954 = N1292 & N1303;
  assign N953 = N1292 & N1304;
  assign N952 = N1293 & N1297;
  assign N951 = N1293 & N1298;
  assign N950 = N1293 & N1299;
  assign N949 = N1293 & N1300;
  assign N948 = N1293 & N1301;
  assign N947 = N1293 & N1302;
  assign N946 = N1293 & N1303;
  assign N945 = N1293 & N1304;
  assign N944 = N1294 & N1297;
  assign N943 = N1294 & N1298;
  assign N942 = N1294 & N1299;
  assign N941 = N1294 & N1300;
  assign N940 = N1294 & N1301;
  assign N939 = N1294 & N1302;
  assign N938 = N1294 & N1303;
  assign N937 = N1294 & N1304;
  assign N936 = N1295 & N1297;
  assign N935 = N1295 & N1298;
  assign N934 = N1295 & N1299;
  assign N933 = N1295 & N1300;
  assign N932 = N1295 & N1301;
  assign N931 = N1295 & N1302;
  assign N930 = N1295 & N1303;
  assign N929 = N1295 & N1304;
  assign N928 = N1296 & N1297;
  assign N927 = N1296 & N1298;
  assign N926 = N1296 & N1299;
  assign N925 = N1296 & N1300;
  assign N924 = N1296 & N1301;
  assign N923 = N1296 & N1302;
  assign N922 = N1296 & N1303;
  assign N921 = N1296 & N1304;
  assign N1319 = yumi_cnt_i[3] & yumi_cnt_i[4];
  assign N1320 = N16 & yumi_cnt_i[4];
  assign N16 = ~yumi_cnt_i[3];
  assign N1321 = yumi_cnt_i[3] & N17;
  assign N17 = ~yumi_cnt_i[4];
  assign N1322 = N18 & N19;
  assign N18 = ~yumi_cnt_i[3];
  assign N19 = ~yumi_cnt_i[4];
  assign N1323 = yumi_cnt_i[5] & N1319;
  assign N1324 = yumi_cnt_i[5] & N1320;
  assign N1325 = yumi_cnt_i[5] & N1321;
  assign N1326 = yumi_cnt_i[5] & N1322;
  assign N1327 = N1255 & N1319;
  assign N1328 = N1255 & N1320;
  assign N1329 = N1255 & N1321;
  assign N1330 = N1255 & N1322;
  assign N1331 = yumi_cnt_i[0] & yumi_cnt_i[1];
  assign N1332 = N20 & yumi_cnt_i[1];
  assign N20 = ~yumi_cnt_i[0];
  assign N1333 = yumi_cnt_i[0] & N21;
  assign N21 = ~yumi_cnt_i[1];
  assign N1334 = N22 & N23;
  assign N22 = ~yumi_cnt_i[0];
  assign N23 = ~yumi_cnt_i[1];
  assign N1335 = yumi_cnt_i[2] & N1331;
  assign N1336 = yumi_cnt_i[2] & N1332;
  assign N1337 = yumi_cnt_i[2] & N1333;
  assign N1338 = yumi_cnt_i[2] & N1334;
  assign N1339 = N1260 & N1331;
  assign N1340 = N1260 & N1332;
  assign N1341 = N1260 & N1333;
  assign N1342 = N1260 & N1334;
  assign N1343 = N1323 & N1336;
  assign N1344 = N1323 & N1337;
  assign N1345 = N1323 & N1338;
  assign N1346 = N1323 & N1342;
  assign N1347 = N1324 & N1335;
  assign N1348 = N1324 & N1336;
  assign N1349 = N1324 & N1337;
  assign N1350 = N1324 & N1338;
  assign N1351 = N1324 & N1339;
  assign N1352 = N1324 & N1340;
  assign N1353 = N1324 & N1341;
  assign N1354 = N1324 & N1342;
  assign N1355 = N1325 & N1335;
  assign N1356 = N1325 & N1336;
  assign N1357 = N1325 & N1337;
  assign N1358 = N1325 & N1338;
  assign N1359 = N1325 & N1339;
  assign N1360 = N1325 & N1340;
  assign N1361 = N1325 & N1341;
  assign N1362 = N1325 & N1342;
  assign N1363 = N1326 & N1335;
  assign N1364 = N1326 & N1336;
  assign N1365 = N1326 & N1337;
  assign N1366 = N1326 & N1338;
  assign N1367 = N1326 & N1339;
  assign N1368 = N1326 & N1340;
  assign N1369 = N1326 & N1341;
  assign N987 = N1326 & N1342;
  assign N986 = N1327 & N1335;
  assign N985 = N1327 & N1336;
  assign N984 = N1327 & N1337;
  assign N983 = N1327 & N1338;
  assign N982 = N1327 & N1339;
  assign N981 = N1327 & N1340;
  assign N980 = N1327 & N1341;
  assign N979 = N1327 & N1342;
  assign N978 = N1328 & N1335;
  assign N977 = N1328 & N1336;
  assign N976 = N1328 & N1337;
  assign N975 = N1328 & N1338;
  assign N974 = N1328 & N1339;
  assign N973 = N1328 & N1340;
  assign N972 = N1328 & N1341;
  assign N971 = N1328 & N1342;
  assign N970 = N1329 & N1335;
  assign N969 = N1329 & N1336;
  assign N968 = N1329 & N1337;
  assign N967 = N1329 & N1338;
  assign N966 = N1329 & N1339;
  assign N965 = N1329 & N1340;
  assign N964 = N1329 & N1341;
  assign N963 = N1329 & N1342;
  assign N962 = N1330 & N1335;
  assign N961 = N1330 & N1336;
  assign N960 = N1330 & N1337;
  assign N959 = N1330 & N1338;
  assign N958 = N1330 & N1339;
  assign N957 = N1330 & N1340;
  assign N956 = N1330 & N1341;
  assign N955 = N1330 & N1342;
  assign { data_o[0:0], data_o[1:1], data_o[2:2], data_o[3:3], data_o[4:4], data_o[5:5], data_o[6:6], data_o[7:7], data_o[8:8], data_o[9:9], data_o[10:10], data_o[11:11], data_o[12:12], data_o[13:13], data_o[14:14], data_o[15:15] } = (N24)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                          (N473)? { data_r[0:0], data_r[1:1], data_r[2:2], data_r[3:3], data_r[4:4], data_r[5:5], data_r[6:6], data_r[7:7], data_r[8:8], data_r[9:9], data_r[10:10], data_r[11:11], data_r[12:12], data_r[13:13], data_r[14:14], data_r[15:15] } : 1'b0;
  assign N24 = N409;
  assign { data_o[16:16], data_o[17:17], data_o[18:18], data_o[19:19], data_o[20:20], data_o[21:21], data_o[22:22], data_o[23:23], data_o[24:24], data_o[25:25], data_o[26:26], data_o[27:27], data_o[28:28], data_o[29:29], data_o[30:30], data_o[31:31] } = (N25)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                              (N474)? { data_r[16:16], data_r[17:17], data_r[18:18], data_r[19:19], data_r[20:20], data_r[21:21], data_r[22:22], data_r[23:23], data_r[24:24], data_r[25:25], data_r[26:26], data_r[27:27], data_r[28:28], data_r[29:29], data_r[30:30], data_r[31:31] } : 1'b0;
  assign N25 = N410;
  assign { data_o[32:32], data_o[33:33], data_o[34:34], data_o[35:35], data_o[36:36], data_o[37:37], data_o[38:38], data_o[39:39], data_o[40:40], data_o[41:41], data_o[42:42], data_o[43:43], data_o[44:44], data_o[45:45], data_o[46:46], data_o[47:47] } = (N26)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                              (N475)? { data_r[32:32], data_r[33:33], data_r[34:34], data_r[35:35], data_r[36:36], data_r[37:37], data_r[38:38], data_r[39:39], data_r[40:40], data_r[41:41], data_r[42:42], data_r[43:43], data_r[44:44], data_r[45:45], data_r[46:46], data_r[47:47] } : 1'b0;
  assign N26 = N411;
  assign { data_o[48:48], data_o[49:49], data_o[50:50], data_o[51:51], data_o[52:52], data_o[53:53], data_o[54:54], data_o[55:55], data_o[56:56], data_o[57:57], data_o[58:58], data_o[59:59], data_o[60:60], data_o[61:61], data_o[62:62], data_o[63:63] } = (N27)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                              (N476)? { data_r[48:48], data_r[49:49], data_r[50:50], data_r[51:51], data_r[52:52], data_r[53:53], data_r[54:54], data_r[55:55], data_r[56:56], data_r[57:57], data_r[58:58], data_r[59:59], data_r[60:60], data_r[61:61], data_r[62:62], data_r[63:63] } : 1'b0;
  assign N27 = N412;
  assign { data_o[64:64], data_o[65:65], data_o[66:66], data_o[67:67], data_o[68:68], data_o[69:69], data_o[70:70], data_o[71:71], data_o[72:72], data_o[73:73], data_o[74:74], data_o[75:75], data_o[76:76], data_o[77:77], data_o[78:78], data_o[79:79] } = (N28)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                              (N477)? { data_r[64:64], data_r[65:65], data_r[66:66], data_r[67:67], data_r[68:68], data_r[69:69], data_r[70:70], data_r[71:71], data_r[72:72], data_r[73:73], data_r[74:74], data_r[75:75], data_r[76:76], data_r[77:77], data_r[78:78], data_r[79:79] } : 1'b0;
  assign N28 = N413;
  assign { data_o[80:80], data_o[81:81], data_o[82:82], data_o[83:83], data_o[84:84], data_o[85:85], data_o[86:86], data_o[87:87], data_o[88:88], data_o[89:89], data_o[90:90], data_o[91:91], data_o[92:92], data_o[93:93], data_o[94:94], data_o[95:95] } = (N29)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                              (N478)? { data_r[80:80], data_r[81:81], data_r[82:82], data_r[83:83], data_r[84:84], data_r[85:85], data_r[86:86], data_r[87:87], data_r[88:88], data_r[89:89], data_r[90:90], data_r[91:91], data_r[92:92], data_r[93:93], data_r[94:94], data_r[95:95] } : 1'b0;
  assign N29 = N414;
  assign { data_o[96:96], data_o[97:97], data_o[98:98], data_o[99:99], data_o[100:100], data_o[101:101], data_o[102:102], data_o[103:103], data_o[104:104], data_o[105:105], data_o[106:106], data_o[107:107], data_o[108:108], data_o[109:109], data_o[110:110], data_o[111:111] } = (N30)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                      (N479)? { data_r[96:96], data_r[97:97], data_r[98:98], data_r[99:99], data_r[100:100], data_r[101:101], data_r[102:102], data_r[103:103], data_r[104:104], data_r[105:105], data_r[106:106], data_r[107:107], data_r[108:108], data_r[109:109], data_r[110:110], data_r[111:111] } : 1'b0;
  assign N30 = N415;
  assign { data_o[112:112], data_o[113:113], data_o[114:114], data_o[115:115], data_o[116:116], data_o[117:117], data_o[118:118], data_o[119:119], data_o[120:120], data_o[121:121], data_o[122:122], data_o[123:123], data_o[124:124], data_o[125:125], data_o[126:126], data_o[127:127] } = (N31)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N480)? { data_r[112:112], data_r[113:113], data_r[114:114], data_r[115:115], data_r[116:116], data_r[117:117], data_r[118:118], data_r[119:119], data_r[120:120], data_r[121:121], data_r[122:122], data_r[123:123], data_r[124:124], data_r[125:125], data_r[126:126], data_r[127:127] } : 1'b0;
  assign N31 = N416;
  assign { data_o[128:128], data_o[129:129], data_o[130:130], data_o[131:131], data_o[132:132], data_o[133:133], data_o[134:134], data_o[135:135], data_o[136:136], data_o[137:137], data_o[138:138], data_o[139:139], data_o[140:140], data_o[141:141], data_o[142:142], data_o[143:143] } = (N32)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N481)? { data_r[128:128], data_r[129:129], data_r[130:130], data_r[131:131], data_r[132:132], data_r[133:133], data_r[134:134], data_r[135:135], data_r[136:136], data_r[137:137], data_r[138:138], data_r[139:139], data_r[140:140], data_r[141:141], data_r[142:142], data_r[143:143] } : 1'b0;
  assign N32 = N417;
  assign { data_o[144:144], data_o[145:145], data_o[146:146], data_o[147:147], data_o[148:148], data_o[149:149], data_o[150:150], data_o[151:151], data_o[152:152], data_o[153:153], data_o[154:154], data_o[155:155], data_o[156:156], data_o[157:157], data_o[158:158], data_o[159:159] } = (N33)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N482)? { data_r[144:144], data_r[145:145], data_r[146:146], data_r[147:147], data_r[148:148], data_r[149:149], data_r[150:150], data_r[151:151], data_r[152:152], data_r[153:153], data_r[154:154], data_r[155:155], data_r[156:156], data_r[157:157], data_r[158:158], data_r[159:159] } : 1'b0;
  assign N33 = N418;
  assign { data_o[160:160], data_o[161:161], data_o[162:162], data_o[163:163], data_o[164:164], data_o[165:165], data_o[166:166], data_o[167:167], data_o[168:168], data_o[169:169], data_o[170:170], data_o[171:171], data_o[172:172], data_o[173:173], data_o[174:174], data_o[175:175] } = (N34)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N483)? { data_r[160:160], data_r[161:161], data_r[162:162], data_r[163:163], data_r[164:164], data_r[165:165], data_r[166:166], data_r[167:167], data_r[168:168], data_r[169:169], data_r[170:170], data_r[171:171], data_r[172:172], data_r[173:173], data_r[174:174], data_r[175:175] } : 1'b0;
  assign N34 = N419;
  assign { data_o[176:176], data_o[177:177], data_o[178:178], data_o[179:179], data_o[180:180], data_o[181:181], data_o[182:182], data_o[183:183], data_o[184:184], data_o[185:185], data_o[186:186], data_o[187:187], data_o[188:188], data_o[189:189], data_o[190:190], data_o[191:191] } = (N35)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N484)? { data_r[176:176], data_r[177:177], data_r[178:178], data_r[179:179], data_r[180:180], data_r[181:181], data_r[182:182], data_r[183:183], data_r[184:184], data_r[185:185], data_r[186:186], data_r[187:187], data_r[188:188], data_r[189:189], data_r[190:190], data_r[191:191] } : 1'b0;
  assign N35 = N420;
  assign { data_o[192:192], data_o[193:193], data_o[194:194], data_o[195:195], data_o[196:196], data_o[197:197], data_o[198:198], data_o[199:199], data_o[200:200], data_o[201:201], data_o[202:202], data_o[203:203], data_o[204:204], data_o[205:205], data_o[206:206], data_o[207:207] } = (N36)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N485)? { data_r[192:192], data_r[193:193], data_r[194:194], data_r[195:195], data_r[196:196], data_r[197:197], data_r[198:198], data_r[199:199], data_r[200:200], data_r[201:201], data_r[202:202], data_r[203:203], data_r[204:204], data_r[205:205], data_r[206:206], data_r[207:207] } : 1'b0;
  assign N36 = N421;
  assign { data_o[208:208], data_o[209:209], data_o[210:210], data_o[211:211], data_o[212:212], data_o[213:213], data_o[214:214], data_o[215:215], data_o[216:216], data_o[217:217], data_o[218:218], data_o[219:219], data_o[220:220], data_o[221:221], data_o[222:222], data_o[223:223] } = (N37)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N486)? { data_r[208:208], data_r[209:209], data_r[210:210], data_r[211:211], data_r[212:212], data_r[213:213], data_r[214:214], data_r[215:215], data_r[216:216], data_r[217:217], data_r[218:218], data_r[219:219], data_r[220:220], data_r[221:221], data_r[222:222], data_r[223:223] } : 1'b0;
  assign N37 = N422;
  assign { data_o[224:224], data_o[225:225], data_o[226:226], data_o[227:227], data_o[228:228], data_o[229:229], data_o[230:230], data_o[231:231], data_o[232:232], data_o[233:233], data_o[234:234], data_o[235:235], data_o[236:236], data_o[237:237], data_o[238:238], data_o[239:239] } = (N38)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N487)? { data_r[224:224], data_r[225:225], data_r[226:226], data_r[227:227], data_r[228:228], data_r[229:229], data_r[230:230], data_r[231:231], data_r[232:232], data_r[233:233], data_r[234:234], data_r[235:235], data_r[236:236], data_r[237:237], data_r[238:238], data_r[239:239] } : 1'b0;
  assign N38 = N423;
  assign { data_o[240:240], data_o[241:241], data_o[242:242], data_o[243:243], data_o[244:244], data_o[245:245], data_o[246:246], data_o[247:247], data_o[248:248], data_o[249:249], data_o[250:250], data_o[251:251], data_o[252:252], data_o[253:253], data_o[254:254], data_o[255:255] } = (N39)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N488)? { data_r[240:240], data_r[241:241], data_r[242:242], data_r[243:243], data_r[244:244], data_r[245:245], data_r[246:246], data_r[247:247], data_r[248:248], data_r[249:249], data_r[250:250], data_r[251:251], data_r[252:252], data_r[253:253], data_r[254:254], data_r[255:255] } : 1'b0;
  assign N39 = N424;
  assign { data_o[256:256], data_o[257:257], data_o[258:258], data_o[259:259], data_o[260:260], data_o[261:261], data_o[262:262], data_o[263:263], data_o[264:264], data_o[265:265], data_o[266:266], data_o[267:267], data_o[268:268], data_o[269:269], data_o[270:270], data_o[271:271] } = (N40)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N489)? { data_r[256:256], data_r[257:257], data_r[258:258], data_r[259:259], data_r[260:260], data_r[261:261], data_r[262:262], data_r[263:263], data_r[264:264], data_r[265:265], data_r[266:266], data_r[267:267], data_r[268:268], data_r[269:269], data_r[270:270], data_r[271:271] } : 1'b0;
  assign N40 = N425;
  assign { data_o[272:272], data_o[273:273], data_o[274:274], data_o[275:275], data_o[276:276], data_o[277:277], data_o[278:278], data_o[279:279], data_o[280:280], data_o[281:281], data_o[282:282], data_o[283:283], data_o[284:284], data_o[285:285], data_o[286:286], data_o[287:287] } = (N41)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N490)? { data_r[272:272], data_r[273:273], data_r[274:274], data_r[275:275], data_r[276:276], data_r[277:277], data_r[278:278], data_r[279:279], data_r[280:280], data_r[281:281], data_r[282:282], data_r[283:283], data_r[284:284], data_r[285:285], data_r[286:286], data_r[287:287] } : 1'b0;
  assign N41 = N426;
  assign { data_o[288:288], data_o[289:289], data_o[290:290], data_o[291:291], data_o[292:292], data_o[293:293], data_o[294:294], data_o[295:295], data_o[296:296], data_o[297:297], data_o[298:298], data_o[299:299], data_o[300:300], data_o[301:301], data_o[302:302], data_o[303:303] } = (N42)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N491)? { data_r[288:288], data_r[289:289], data_r[290:290], data_r[291:291], data_r[292:292], data_r[293:293], data_r[294:294], data_r[295:295], data_r[296:296], data_r[297:297], data_r[298:298], data_r[299:299], data_r[300:300], data_r[301:301], data_r[302:302], data_r[303:303] } : 1'b0;
  assign N42 = N427;
  assign { data_o[304:304], data_o[305:305], data_o[306:306], data_o[307:307], data_o[308:308], data_o[309:309], data_o[310:310], data_o[311:311], data_o[312:312], data_o[313:313], data_o[314:314], data_o[315:315], data_o[316:316], data_o[317:317], data_o[318:318], data_o[319:319] } = (N43)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N492)? { data_r[304:304], data_r[305:305], data_r[306:306], data_r[307:307], data_r[308:308], data_r[309:309], data_r[310:310], data_r[311:311], data_r[312:312], data_r[313:313], data_r[314:314], data_r[315:315], data_r[316:316], data_r[317:317], data_r[318:318], data_r[319:319] } : 1'b0;
  assign N43 = N428;
  assign { data_o[320:320], data_o[321:321], data_o[322:322], data_o[323:323], data_o[324:324], data_o[325:325], data_o[326:326], data_o[327:327], data_o[328:328], data_o[329:329], data_o[330:330], data_o[331:331], data_o[332:332], data_o[333:333], data_o[334:334], data_o[335:335] } = (N44)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N493)? { data_r[320:320], data_r[321:321], data_r[322:322], data_r[323:323], data_r[324:324], data_r[325:325], data_r[326:326], data_r[327:327], data_r[328:328], data_r[329:329], data_r[330:330], data_r[331:331], data_r[332:332], data_r[333:333], data_r[334:334], data_r[335:335] } : 1'b0;
  assign N44 = N429;
  assign { data_o[336:336], data_o[337:337], data_o[338:338], data_o[339:339], data_o[340:340], data_o[341:341], data_o[342:342], data_o[343:343], data_o[344:344], data_o[345:345], data_o[346:346], data_o[347:347], data_o[348:348], data_o[349:349], data_o[350:350], data_o[351:351] } = (N45)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N494)? { data_r[336:336], data_r[337:337], data_r[338:338], data_r[339:339], data_r[340:340], data_r[341:341], data_r[342:342], data_r[343:343], data_r[344:344], data_r[345:345], data_r[346:346], data_r[347:347], data_r[348:348], data_r[349:349], data_r[350:350], data_r[351:351] } : 1'b0;
  assign N45 = N430;
  assign { data_o[352:352], data_o[353:353], data_o[354:354], data_o[355:355], data_o[356:356], data_o[357:357], data_o[358:358], data_o[359:359], data_o[360:360], data_o[361:361], data_o[362:362], data_o[363:363], data_o[364:364], data_o[365:365], data_o[366:366], data_o[367:367] } = (N46)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N495)? { data_r[352:352], data_r[353:353], data_r[354:354], data_r[355:355], data_r[356:356], data_r[357:357], data_r[358:358], data_r[359:359], data_r[360:360], data_r[361:361], data_r[362:362], data_r[363:363], data_r[364:364], data_r[365:365], data_r[366:366], data_r[367:367] } : 1'b0;
  assign N46 = N431;
  assign { data_o[368:368], data_o[369:369], data_o[370:370], data_o[371:371], data_o[372:372], data_o[373:373], data_o[374:374], data_o[375:375], data_o[376:376], data_o[377:377], data_o[378:378], data_o[379:379], data_o[380:380], data_o[381:381], data_o[382:382], data_o[383:383] } = (N47)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N496)? { data_r[368:368], data_r[369:369], data_r[370:370], data_r[371:371], data_r[372:372], data_r[373:373], data_r[374:374], data_r[375:375], data_r[376:376], data_r[377:377], data_r[378:378], data_r[379:379], data_r[380:380], data_r[381:381], data_r[382:382], data_r[383:383] } : 1'b0;
  assign N47 = N432;
  assign { data_o[384:384], data_o[385:385], data_o[386:386], data_o[387:387], data_o[388:388], data_o[389:389], data_o[390:390], data_o[391:391], data_o[392:392], data_o[393:393], data_o[394:394], data_o[395:395], data_o[396:396], data_o[397:397], data_o[398:398], data_o[399:399] } = (N48)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N497)? { data_r[384:384], data_r[385:385], data_r[386:386], data_r[387:387], data_r[388:388], data_r[389:389], data_r[390:390], data_r[391:391], data_r[392:392], data_r[393:393], data_r[394:394], data_r[395:395], data_r[396:396], data_r[397:397], data_r[398:398], data_r[399:399] } : 1'b0;
  assign N48 = N433;
  assign { data_o[400:400], data_o[401:401], data_o[402:402], data_o[403:403], data_o[404:404], data_o[405:405], data_o[406:406], data_o[407:407], data_o[408:408], data_o[409:409], data_o[410:410], data_o[411:411], data_o[412:412], data_o[413:413], data_o[414:414], data_o[415:415] } = (N49)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N498)? { data_r[400:400], data_r[401:401], data_r[402:402], data_r[403:403], data_r[404:404], data_r[405:405], data_r[406:406], data_r[407:407], data_r[408:408], data_r[409:409], data_r[410:410], data_r[411:411], data_r[412:412], data_r[413:413], data_r[414:414], data_r[415:415] } : 1'b0;
  assign N49 = N434;
  assign { data_o[416:416], data_o[417:417], data_o[418:418], data_o[419:419], data_o[420:420], data_o[421:421], data_o[422:422], data_o[423:423], data_o[424:424], data_o[425:425], data_o[426:426], data_o[427:427], data_o[428:428], data_o[429:429], data_o[430:430], data_o[431:431] } = (N50)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N499)? { data_r[416:416], data_r[417:417], data_r[418:418], data_r[419:419], data_r[420:420], data_r[421:421], data_r[422:422], data_r[423:423], data_r[424:424], data_r[425:425], data_r[426:426], data_r[427:427], data_r[428:428], data_r[429:429], data_r[430:430], data_r[431:431] } : 1'b0;
  assign N50 = N435;
  assign { data_o[432:432], data_o[433:433], data_o[434:434], data_o[435:435], data_o[436:436], data_o[437:437], data_o[438:438], data_o[439:439], data_o[440:440], data_o[441:441], data_o[442:442], data_o[443:443], data_o[444:444], data_o[445:445], data_o[446:446], data_o[447:447] } = (N51)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N500)? { data_r[432:432], data_r[433:433], data_r[434:434], data_r[435:435], data_r[436:436], data_r[437:437], data_r[438:438], data_r[439:439], data_r[440:440], data_r[441:441], data_r[442:442], data_r[443:443], data_r[444:444], data_r[445:445], data_r[446:446], data_r[447:447] } : 1'b0;
  assign N51 = N436;
  assign { data_o[448:448], data_o[449:449], data_o[450:450], data_o[451:451], data_o[452:452], data_o[453:453], data_o[454:454], data_o[455:455], data_o[456:456], data_o[457:457], data_o[458:458], data_o[459:459], data_o[460:460], data_o[461:461], data_o[462:462], data_o[463:463] } = (N52)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N501)? { data_r[448:448], data_r[449:449], data_r[450:450], data_r[451:451], data_r[452:452], data_r[453:453], data_r[454:454], data_r[455:455], data_r[456:456], data_r[457:457], data_r[458:458], data_r[459:459], data_r[460:460], data_r[461:461], data_r[462:462], data_r[463:463] } : 1'b0;
  assign N52 = N437;
  assign { data_o[464:464], data_o[465:465], data_o[466:466], data_o[467:467], data_o[468:468], data_o[469:469], data_o[470:470], data_o[471:471], data_o[472:472], data_o[473:473], data_o[474:474], data_o[475:475], data_o[476:476], data_o[477:477], data_o[478:478], data_o[479:479] } = (N53)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N502)? { data_r[464:464], data_r[465:465], data_r[466:466], data_r[467:467], data_r[468:468], data_r[469:469], data_r[470:470], data_r[471:471], data_r[472:472], data_r[473:473], data_r[474:474], data_r[475:475], data_r[476:476], data_r[477:477], data_r[478:478], data_r[479:479] } : 1'b0;
  assign N53 = N438;
  assign { data_o[480:480], data_o[481:481], data_o[482:482], data_o[483:483], data_o[484:484], data_o[485:485], data_o[486:486], data_o[487:487], data_o[488:488], data_o[489:489], data_o[490:490], data_o[491:491], data_o[492:492], data_o[493:493], data_o[494:494], data_o[495:495] } = (N54)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N503)? { data_r[480:480], data_r[481:481], data_r[482:482], data_r[483:483], data_r[484:484], data_r[485:485], data_r[486:486], data_r[487:487], data_r[488:488], data_r[489:489], data_r[490:490], data_r[491:491], data_r[492:492], data_r[493:493], data_r[494:494], data_r[495:495] } : 1'b0;
  assign N54 = N439;
  assign { data_o[496:496], data_o[497:497], data_o[498:498], data_o[499:499], data_o[500:500], data_o[501:501], data_o[502:502], data_o[503:503], data_o[504:504], data_o[505:505], data_o[506:506], data_o[507:507], data_o[508:508], data_o[509:509], data_o[510:510], data_o[511:511] } = (N55)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                                              (N504)? { data_r[496:496], data_r[497:497], data_r[498:498], data_r[499:499], data_r[500:500], data_r[501:501], data_r[502:502], data_r[503:503], data_r[504:504], data_r[505:505], data_r[506:506], data_r[507:507], data_r[508:508], data_r[509:509], data_r[510:510], data_r[511:511] } : 1'b0;
  assign N55 = N440;
  assign { data_n_32__0_, data_n_32__1_, data_n_32__2_, data_n_32__3_, data_n_32__4_, data_n_32__5_, data_n_32__6_, data_n_32__7_, data_n_32__8_, data_n_32__9_, data_n_32__10_, data_n_32__11_, data_n_32__12_, data_n_32__13_, data_n_32__14_, data_n_32__15_ } = (N56)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N505)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N56 = N441;
  assign { data_n_33__0_, data_n_33__1_, data_n_33__2_, data_n_33__3_, data_n_33__4_, data_n_33__5_, data_n_33__6_, data_n_33__7_, data_n_33__8_, data_n_33__9_, data_n_33__10_, data_n_33__11_, data_n_33__12_, data_n_33__13_, data_n_33__14_, data_n_33__15_ } = (N57)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N506)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N57 = N442;
  assign { data_n_34__0_, data_n_34__1_, data_n_34__2_, data_n_34__3_, data_n_34__4_, data_n_34__5_, data_n_34__6_, data_n_34__7_, data_n_34__8_, data_n_34__9_, data_n_34__10_, data_n_34__11_, data_n_34__12_, data_n_34__13_, data_n_34__14_, data_n_34__15_ } = (N58)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N507)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N58 = N443;
  assign { data_n_35__0_, data_n_35__1_, data_n_35__2_, data_n_35__3_, data_n_35__4_, data_n_35__5_, data_n_35__6_, data_n_35__7_, data_n_35__8_, data_n_35__9_, data_n_35__10_, data_n_35__11_, data_n_35__12_, data_n_35__13_, data_n_35__14_, data_n_35__15_ } = (N59)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N508)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N59 = N444;
  assign { data_n_36__0_, data_n_36__1_, data_n_36__2_, data_n_36__3_, data_n_36__4_, data_n_36__5_, data_n_36__6_, data_n_36__7_, data_n_36__8_, data_n_36__9_, data_n_36__10_, data_n_36__11_, data_n_36__12_, data_n_36__13_, data_n_36__14_, data_n_36__15_ } = (N60)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N509)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N60 = N445;
  assign { data_n_37__0_, data_n_37__1_, data_n_37__2_, data_n_37__3_, data_n_37__4_, data_n_37__5_, data_n_37__6_, data_n_37__7_, data_n_37__8_, data_n_37__9_, data_n_37__10_, data_n_37__11_, data_n_37__12_, data_n_37__13_, data_n_37__14_, data_n_37__15_ } = (N61)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N510)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N61 = N446;
  assign { data_n_38__0_, data_n_38__1_, data_n_38__2_, data_n_38__3_, data_n_38__4_, data_n_38__5_, data_n_38__6_, data_n_38__7_, data_n_38__8_, data_n_38__9_, data_n_38__10_, data_n_38__11_, data_n_38__12_, data_n_38__13_, data_n_38__14_, data_n_38__15_ } = (N62)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N511)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N62 = N447;
  assign { data_n_39__0_, data_n_39__1_, data_n_39__2_, data_n_39__3_, data_n_39__4_, data_n_39__5_, data_n_39__6_, data_n_39__7_, data_n_39__8_, data_n_39__9_, data_n_39__10_, data_n_39__11_, data_n_39__12_, data_n_39__13_, data_n_39__14_, data_n_39__15_ } = (N63)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N512)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N63 = N448;
  assign { data_n_40__0_, data_n_40__1_, data_n_40__2_, data_n_40__3_, data_n_40__4_, data_n_40__5_, data_n_40__6_, data_n_40__7_, data_n_40__8_, data_n_40__9_, data_n_40__10_, data_n_40__11_, data_n_40__12_, data_n_40__13_, data_n_40__14_, data_n_40__15_ } = (N64)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N513)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N64 = N449;
  assign { data_n_41__0_, data_n_41__1_, data_n_41__2_, data_n_41__3_, data_n_41__4_, data_n_41__5_, data_n_41__6_, data_n_41__7_, data_n_41__8_, data_n_41__9_, data_n_41__10_, data_n_41__11_, data_n_41__12_, data_n_41__13_, data_n_41__14_, data_n_41__15_ } = (N65)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N514)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N65 = N450;
  assign { data_n_42__0_, data_n_42__1_, data_n_42__2_, data_n_42__3_, data_n_42__4_, data_n_42__5_, data_n_42__6_, data_n_42__7_, data_n_42__8_, data_n_42__9_, data_n_42__10_, data_n_42__11_, data_n_42__12_, data_n_42__13_, data_n_42__14_, data_n_42__15_ } = (N66)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N515)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N66 = N451;
  assign { data_n_43__0_, data_n_43__1_, data_n_43__2_, data_n_43__3_, data_n_43__4_, data_n_43__5_, data_n_43__6_, data_n_43__7_, data_n_43__8_, data_n_43__9_, data_n_43__10_, data_n_43__11_, data_n_43__12_, data_n_43__13_, data_n_43__14_, data_n_43__15_ } = (N67)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N516)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N67 = N452;
  assign { data_n_44__0_, data_n_44__1_, data_n_44__2_, data_n_44__3_, data_n_44__4_, data_n_44__5_, data_n_44__6_, data_n_44__7_, data_n_44__8_, data_n_44__9_, data_n_44__10_, data_n_44__11_, data_n_44__12_, data_n_44__13_, data_n_44__14_, data_n_44__15_ } = (N68)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N517)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N68 = N453;
  assign { data_n_45__0_, data_n_45__1_, data_n_45__2_, data_n_45__3_, data_n_45__4_, data_n_45__5_, data_n_45__6_, data_n_45__7_, data_n_45__8_, data_n_45__9_, data_n_45__10_, data_n_45__11_, data_n_45__12_, data_n_45__13_, data_n_45__14_, data_n_45__15_ } = (N69)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N518)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N69 = N454;
  assign { data_n_46__0_, data_n_46__1_, data_n_46__2_, data_n_46__3_, data_n_46__4_, data_n_46__5_, data_n_46__6_, data_n_46__7_, data_n_46__8_, data_n_46__9_, data_n_46__10_, data_n_46__11_, data_n_46__12_, data_n_46__13_, data_n_46__14_, data_n_46__15_ } = (N70)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N519)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N70 = N455;
  assign { data_n_47__0_, data_n_47__1_, data_n_47__2_, data_n_47__3_, data_n_47__4_, data_n_47__5_, data_n_47__6_, data_n_47__7_, data_n_47__8_, data_n_47__9_, data_n_47__10_, data_n_47__11_, data_n_47__12_, data_n_47__13_, data_n_47__14_, data_n_47__15_ } = (N71)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N520)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N71 = N456;
  assign { data_n_48__0_, data_n_48__1_, data_n_48__2_, data_n_48__3_, data_n_48__4_, data_n_48__5_, data_n_48__6_, data_n_48__7_, data_n_48__8_, data_n_48__9_, data_n_48__10_, data_n_48__11_, data_n_48__12_, data_n_48__13_, data_n_48__14_, data_n_48__15_ } = (N72)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N521)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N72 = N457;
  assign { data_n_49__0_, data_n_49__1_, data_n_49__2_, data_n_49__3_, data_n_49__4_, data_n_49__5_, data_n_49__6_, data_n_49__7_, data_n_49__8_, data_n_49__9_, data_n_49__10_, data_n_49__11_, data_n_49__12_, data_n_49__13_, data_n_49__14_, data_n_49__15_ } = (N73)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N522)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N73 = N458;
  assign { data_n_50__0_, data_n_50__1_, data_n_50__2_, data_n_50__3_, data_n_50__4_, data_n_50__5_, data_n_50__6_, data_n_50__7_, data_n_50__8_, data_n_50__9_, data_n_50__10_, data_n_50__11_, data_n_50__12_, data_n_50__13_, data_n_50__14_, data_n_50__15_ } = (N74)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N523)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N74 = N459;
  assign { data_n_51__0_, data_n_51__1_, data_n_51__2_, data_n_51__3_, data_n_51__4_, data_n_51__5_, data_n_51__6_, data_n_51__7_, data_n_51__8_, data_n_51__9_, data_n_51__10_, data_n_51__11_, data_n_51__12_, data_n_51__13_, data_n_51__14_, data_n_51__15_ } = (N75)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N524)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N75 = N460;
  assign { data_n_52__0_, data_n_52__1_, data_n_52__2_, data_n_52__3_, data_n_52__4_, data_n_52__5_, data_n_52__6_, data_n_52__7_, data_n_52__8_, data_n_52__9_, data_n_52__10_, data_n_52__11_, data_n_52__12_, data_n_52__13_, data_n_52__14_, data_n_52__15_ } = (N76)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N525)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N76 = N461;
  assign { data_n_53__0_, data_n_53__1_, data_n_53__2_, data_n_53__3_, data_n_53__4_, data_n_53__5_, data_n_53__6_, data_n_53__7_, data_n_53__8_, data_n_53__9_, data_n_53__10_, data_n_53__11_, data_n_53__12_, data_n_53__13_, data_n_53__14_, data_n_53__15_ } = (N77)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N526)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N77 = N462;
  assign { data_n_54__0_, data_n_54__1_, data_n_54__2_, data_n_54__3_, data_n_54__4_, data_n_54__5_, data_n_54__6_, data_n_54__7_, data_n_54__8_, data_n_54__9_, data_n_54__10_, data_n_54__11_, data_n_54__12_, data_n_54__13_, data_n_54__14_, data_n_54__15_ } = (N78)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N527)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N78 = N463;
  assign { data_n_55__0_, data_n_55__1_, data_n_55__2_, data_n_55__3_, data_n_55__4_, data_n_55__5_, data_n_55__6_, data_n_55__7_, data_n_55__8_, data_n_55__9_, data_n_55__10_, data_n_55__11_, data_n_55__12_, data_n_55__13_, data_n_55__14_, data_n_55__15_ } = (N79)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N528)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N79 = N464;
  assign { data_n_56__0_, data_n_56__1_, data_n_56__2_, data_n_56__3_, data_n_56__4_, data_n_56__5_, data_n_56__6_, data_n_56__7_, data_n_56__8_, data_n_56__9_, data_n_56__10_, data_n_56__11_, data_n_56__12_, data_n_56__13_, data_n_56__14_, data_n_56__15_ } = (N80)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N529)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N80 = N465;
  assign { data_n_57__0_, data_n_57__1_, data_n_57__2_, data_n_57__3_, data_n_57__4_, data_n_57__5_, data_n_57__6_, data_n_57__7_, data_n_57__8_, data_n_57__9_, data_n_57__10_, data_n_57__11_, data_n_57__12_, data_n_57__13_, data_n_57__14_, data_n_57__15_ } = (N81)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N530)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N81 = N466;
  assign { data_n_58__0_, data_n_58__1_, data_n_58__2_, data_n_58__3_, data_n_58__4_, data_n_58__5_, data_n_58__6_, data_n_58__7_, data_n_58__8_, data_n_58__9_, data_n_58__10_, data_n_58__11_, data_n_58__12_, data_n_58__13_, data_n_58__14_, data_n_58__15_ } = (N82)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N531)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N82 = N467;
  assign { data_n_59__0_, data_n_59__1_, data_n_59__2_, data_n_59__3_, data_n_59__4_, data_n_59__5_, data_n_59__6_, data_n_59__7_, data_n_59__8_, data_n_59__9_, data_n_59__10_, data_n_59__11_, data_n_59__12_, data_n_59__13_, data_n_59__14_, data_n_59__15_ } = (N83)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N532)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N83 = N468;
  assign { data_n_60__0_, data_n_60__1_, data_n_60__2_, data_n_60__3_, data_n_60__4_, data_n_60__5_, data_n_60__6_, data_n_60__7_, data_n_60__8_, data_n_60__9_, data_n_60__10_, data_n_60__11_, data_n_60__12_, data_n_60__13_, data_n_60__14_, data_n_60__15_ } = (N84)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N533)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N84 = N469;
  assign { data_n_61__0_, data_n_61__1_, data_n_61__2_, data_n_61__3_, data_n_61__4_, data_n_61__5_, data_n_61__6_, data_n_61__7_, data_n_61__8_, data_n_61__9_, data_n_61__10_, data_n_61__11_, data_n_61__12_, data_n_61__13_, data_n_61__14_, data_n_61__15_ } = (N85)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N534)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N85 = N470;
  assign { data_n_62__0_, data_n_62__1_, data_n_62__2_, data_n_62__3_, data_n_62__4_, data_n_62__5_, data_n_62__6_, data_n_62__7_, data_n_62__8_, data_n_62__9_, data_n_62__10_, data_n_62__11_, data_n_62__12_, data_n_62__13_, data_n_62__14_, data_n_62__15_ } = (N86)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N535)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N86 = N471;
  assign { data_n_63__0_, data_n_63__1_, data_n_63__2_, data_n_63__3_, data_n_63__4_, data_n_63__5_, data_n_63__6_, data_n_63__7_, data_n_63__8_, data_n_63__9_, data_n_63__10_, data_n_63__11_, data_n_63__12_, data_n_63__13_, data_n_63__14_, data_n_63__15_ } = (N87)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15] } : 
                                                                                                                                                                                                                                                                    (N536)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N87 = N472;
  assign valid_o[0] = (N88)? N601 : 
                      (N602)? valid_r[0] : 1'b0;
  assign N88 = N537;
  assign valid_o[1] = (N89)? N601 : 
                      (N603)? valid_r[1] : 1'b0;
  assign N89 = N538;
  assign valid_o[2] = (N90)? N601 : 
                      (N604)? valid_r[2] : 1'b0;
  assign N90 = N539;
  assign valid_o[3] = (N91)? N601 : 
                      (N605)? valid_r[3] : 1'b0;
  assign N91 = N540;
  assign valid_o[4] = (N92)? N601 : 
                      (N606)? valid_r[4] : 1'b0;
  assign N92 = N541;
  assign valid_o[5] = (N93)? N601 : 
                      (N607)? valid_r[5] : 1'b0;
  assign N93 = N542;
  assign valid_o[6] = (N94)? N601 : 
                      (N608)? valid_r[6] : 1'b0;
  assign N94 = N543;
  assign valid_o[7] = (N95)? N601 : 
                      (N609)? valid_r[7] : 1'b0;
  assign N95 = N544;
  assign valid_o[8] = (N96)? N601 : 
                      (N610)? valid_r[8] : 1'b0;
  assign N96 = N545;
  assign valid_o[9] = (N97)? N601 : 
                      (N611)? valid_r[9] : 1'b0;
  assign N97 = N546;
  assign valid_o[10] = (N98)? N601 : 
                       (N612)? valid_r[10] : 1'b0;
  assign N98 = N547;
  assign valid_o[11] = (N99)? N601 : 
                       (N613)? valid_r[11] : 1'b0;
  assign N99 = N548;
  assign valid_o[12] = (N100)? N601 : 
                       (N614)? valid_r[12] : 1'b0;
  assign N100 = N549;
  assign valid_o[13] = (N101)? N601 : 
                       (N615)? valid_r[13] : 1'b0;
  assign N101 = N550;
  assign valid_o[14] = (N102)? N601 : 
                       (N616)? valid_r[14] : 1'b0;
  assign N102 = N551;
  assign valid_o[15] = (N103)? N601 : 
                       (N617)? valid_r[15] : 1'b0;
  assign N103 = N552;
  assign valid_o[16] = (N104)? N601 : 
                       (N618)? valid_r[16] : 1'b0;
  assign N104 = N553;
  assign valid_o[17] = (N105)? N601 : 
                       (N619)? valid_r[17] : 1'b0;
  assign N105 = N554;
  assign valid_o[18] = (N106)? N601 : 
                       (N620)? valid_r[18] : 1'b0;
  assign N106 = N555;
  assign valid_o[19] = (N107)? N601 : 
                       (N621)? valid_r[19] : 1'b0;
  assign N107 = N556;
  assign valid_o[20] = (N108)? N601 : 
                       (N622)? valid_r[20] : 1'b0;
  assign N108 = N557;
  assign valid_o[21] = (N109)? N601 : 
                       (N623)? valid_r[21] : 1'b0;
  assign N109 = N558;
  assign valid_o[22] = (N110)? N601 : 
                       (N624)? valid_r[22] : 1'b0;
  assign N110 = N559;
  assign valid_o[23] = (N111)? N601 : 
                       (N625)? valid_r[23] : 1'b0;
  assign N111 = N560;
  assign valid_o[24] = (N112)? N601 : 
                       (N626)? valid_r[24] : 1'b0;
  assign N112 = N561;
  assign valid_o[25] = (N113)? N601 : 
                       (N627)? valid_r[25] : 1'b0;
  assign N113 = N562;
  assign valid_o[26] = (N114)? N601 : 
                       (N628)? valid_r[26] : 1'b0;
  assign N114 = N563;
  assign valid_o[27] = (N115)? N601 : 
                       (N629)? valid_r[27] : 1'b0;
  assign N115 = N564;
  assign valid_o[28] = (N116)? N601 : 
                       (N630)? valid_r[28] : 1'b0;
  assign N116 = N565;
  assign valid_o[29] = (N117)? N601 : 
                       (N631)? valid_r[29] : 1'b0;
  assign N117 = N566;
  assign valid_o[30] = (N118)? N601 : 
                       (N632)? valid_r[30] : 1'b0;
  assign N118 = N567;
  assign valid_o[31] = (N119)? N601 : 
                       (N633)? valid_r[31] : 1'b0;
  assign N119 = N568;
  assign valid_n[32] = (N120)? N601 : 
                       (N634)? 1'b0 : 1'b0;
  assign N120 = N569;
  assign valid_n[33] = (N121)? N601 : 
                       (N635)? 1'b0 : 1'b0;
  assign N121 = N570;
  assign valid_n[34] = (N122)? N601 : 
                       (N636)? 1'b0 : 1'b0;
  assign N122 = N571;
  assign valid_n[35] = (N123)? N601 : 
                       (N637)? 1'b0 : 1'b0;
  assign N123 = N572;
  assign valid_n[36] = (N124)? N601 : 
                       (N638)? 1'b0 : 1'b0;
  assign N124 = N573;
  assign valid_n[37] = (N125)? N601 : 
                       (N639)? 1'b0 : 1'b0;
  assign N125 = N574;
  assign valid_n[38] = (N126)? N601 : 
                       (N640)? 1'b0 : 1'b0;
  assign N126 = N575;
  assign valid_n[39] = (N127)? N601 : 
                       (N641)? 1'b0 : 1'b0;
  assign N127 = N576;
  assign valid_n[40] = (N128)? N601 : 
                       (N642)? 1'b0 : 1'b0;
  assign N128 = N577;
  assign valid_n[41] = (N129)? N601 : 
                       (N643)? 1'b0 : 1'b0;
  assign N129 = N578;
  assign valid_n[42] = (N130)? N601 : 
                       (N644)? 1'b0 : 1'b0;
  assign N130 = N579;
  assign valid_n[43] = (N131)? N601 : 
                       (N645)? 1'b0 : 1'b0;
  assign N131 = N580;
  assign valid_n[44] = (N132)? N601 : 
                       (N646)? 1'b0 : 1'b0;
  assign N132 = N581;
  assign valid_n[45] = (N133)? N601 : 
                       (N647)? 1'b0 : 1'b0;
  assign N133 = N582;
  assign valid_n[46] = (N134)? N601 : 
                       (N648)? 1'b0 : 1'b0;
  assign N134 = N583;
  assign valid_n[47] = (N135)? N601 : 
                       (N649)? 1'b0 : 1'b0;
  assign N135 = N584;
  assign valid_n[48] = (N136)? N601 : 
                       (N650)? 1'b0 : 1'b0;
  assign N136 = N585;
  assign valid_n[49] = (N137)? N601 : 
                       (N651)? 1'b0 : 1'b0;
  assign N137 = N586;
  assign valid_n[50] = (N138)? N601 : 
                       (N652)? 1'b0 : 1'b0;
  assign N138 = N587;
  assign valid_n[51] = (N139)? N601 : 
                       (N653)? 1'b0 : 1'b0;
  assign N139 = N588;
  assign valid_n[52] = (N140)? N601 : 
                       (N654)? 1'b0 : 1'b0;
  assign N140 = N589;
  assign valid_n[53] = (N141)? N601 : 
                       (N655)? 1'b0 : 1'b0;
  assign N141 = N590;
  assign valid_n[54] = (N142)? N601 : 
                       (N656)? 1'b0 : 1'b0;
  assign N142 = N591;
  assign valid_n[55] = (N143)? N601 : 
                       (N657)? 1'b0 : 1'b0;
  assign N143 = N592;
  assign valid_n[56] = (N144)? N601 : 
                       (N658)? 1'b0 : 1'b0;
  assign N144 = N593;
  assign valid_n[57] = (N145)? N601 : 
                       (N659)? 1'b0 : 1'b0;
  assign N145 = N594;
  assign valid_n[58] = (N146)? N601 : 
                       (N660)? 1'b0 : 1'b0;
  assign N146 = N595;
  assign valid_n[59] = (N147)? N601 : 
                       (N661)? 1'b0 : 1'b0;
  assign N147 = N596;
  assign valid_n[60] = (N148)? N601 : 
                       (N662)? 1'b0 : 1'b0;
  assign N148 = N597;
  assign valid_n[61] = (N149)? N601 : 
                       (N663)? 1'b0 : 1'b0;
  assign N149 = N598;
  assign valid_n[62] = (N150)? N601 : 
                       (N664)? 1'b0 : 1'b0;
  assign N150 = N599;
  assign valid_n[63] = (N151)? N601 : 
                       (N665)? 1'b0 : 1'b0;
  assign N151 = N600;
  assign data_nn[31:16] = (N152)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                          (N153)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                          (N154)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                          (N155)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                          (N156)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                          (N157)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                          (N158)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                          (N159)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                          (N160)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                          (N161)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                          (N162)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                          (N163)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                          (N164)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                          (N165)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                          (N166)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                          (N167)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                          (N168)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                          (N169)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                          (N170)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                          (N171)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                          (N172)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                          (N173)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                          (N174)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                          (N175)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                          (N176)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                          (N177)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                          (N178)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                          (N179)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                          (N180)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                          (N181)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                          (N182)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                          (N183)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                          (N184)? data_o[511:496] : 
                          (N185)? data_o[495:480] : 
                          (N186)? data_o[479:464] : 
                          (N187)? data_o[463:448] : 
                          (N188)? data_o[447:432] : 
                          (N189)? data_o[431:416] : 
                          (N190)? data_o[415:400] : 
                          (N191)? data_o[399:384] : 
                          (N192)? data_o[383:368] : 
                          (N193)? data_o[367:352] : 
                          (N194)? data_o[351:336] : 
                          (N195)? data_o[335:320] : 
                          (N196)? data_o[319:304] : 
                          (N197)? data_o[303:288] : 
                          (N198)? data_o[287:272] : 
                          (N199)? data_o[271:256] : 
                          (N200)? data_o[255:240] : 
                          (N201)? data_o[239:224] : 
                          (N202)? data_o[223:208] : 
                          (N203)? data_o[207:192] : 
                          (N204)? data_o[191:176] : 
                          (N205)? data_o[175:160] : 
                          (N206)? data_o[159:144] : 
                          (N207)? data_o[143:128] : 
                          (N208)? data_o[127:112] : 
                          (N209)? data_o[111:96] : 
                          (N210)? data_o[95:80] : 
                          (N211)? data_o[79:64] : 
                          (N212)? data_o[63:48] : 
                          (N213)? data_o[47:32] : 
                          (N214)? data_o[31:16] : 1'b0;
  assign N152 = N1343;
  assign N153 = N1344;
  assign N154 = N1345;
  assign N155 = N1265;
  assign N156 = N1266;
  assign N157 = N841;
  assign N158 = N840;
  assign N159 = N1347;
  assign N160 = N1348;
  assign N161 = N1349;
  assign N162 = N1350;
  assign N163 = N839;
  assign N164 = N838;
  assign N165 = N837;
  assign N166 = N836;
  assign N167 = N1355;
  assign N168 = N1356;
  assign N169 = N1357;
  assign N170 = N1358;
  assign N171 = N835;
  assign N172 = N834;
  assign N173 = N833;
  assign N174 = N832;
  assign N175 = N1363;
  assign N176 = N1364;
  assign N177 = N1365;
  assign N178 = N1366;
  assign N179 = N831;
  assign N180 = N830;
  assign N181 = N829;
  assign N182 = N828;
  assign N183 = N827;
  assign N184 = N826;
  assign N185 = N825;
  assign N186 = N824;
  assign N187 = N823;
  assign N188 = N822;
  assign N189 = N821;
  assign N190 = N820;
  assign N191 = N819;
  assign N192 = N818;
  assign N193 = N817;
  assign N194 = N816;
  assign N195 = N815;
  assign N196 = N814;
  assign N197 = N813;
  assign N198 = N812;
  assign N199 = N811;
  assign N200 = N810;
  assign N201 = N809;
  assign N202 = N808;
  assign N203 = N807;
  assign N204 = N806;
  assign N205 = N805;
  assign N206 = N804;
  assign N207 = N803;
  assign N208 = N802;
  assign N209 = N801;
  assign N210 = N800;
  assign N211 = N799;
  assign N212 = N798;
  assign N213 = N797;
  assign N214 = N796;
  assign data_nn[47:32] = (N153)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                          (N154)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                          (N155)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                          (N156)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                          (N157)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                          (N158)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                          (N159)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                          (N160)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                          (N161)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                          (N162)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                          (N163)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                          (N164)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                          (N165)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                          (N166)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                          (N167)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                          (N168)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                          (N169)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                          (N170)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                          (N171)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                          (N172)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                          (N173)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                          (N174)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                          (N175)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                          (N176)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                          (N177)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                          (N178)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                          (N179)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                          (N180)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                          (N181)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                          (N182)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                          (N183)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                          (N184)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                          (N185)? data_o[511:496] : 
                          (N186)? data_o[495:480] : 
                          (N187)? data_o[479:464] : 
                          (N188)? data_o[463:448] : 
                          (N189)? data_o[447:432] : 
                          (N190)? data_o[431:416] : 
                          (N191)? data_o[415:400] : 
                          (N192)? data_o[399:384] : 
                          (N193)? data_o[383:368] : 
                          (N194)? data_o[367:352] : 
                          (N195)? data_o[351:336] : 
                          (N196)? data_o[335:320] : 
                          (N197)? data_o[319:304] : 
                          (N198)? data_o[303:288] : 
                          (N199)? data_o[287:272] : 
                          (N200)? data_o[271:256] : 
                          (N201)? data_o[255:240] : 
                          (N202)? data_o[239:224] : 
                          (N203)? data_o[223:208] : 
                          (N204)? data_o[207:192] : 
                          (N205)? data_o[191:176] : 
                          (N206)? data_o[175:160] : 
                          (N207)? data_o[159:144] : 
                          (N208)? data_o[143:128] : 
                          (N209)? data_o[127:112] : 
                          (N210)? data_o[111:96] : 
                          (N211)? data_o[95:80] : 
                          (N212)? data_o[79:64] : 
                          (N213)? data_o[63:48] : 
                          (N214)? data_o[47:32] : 1'b0;
  assign data_nn[63:48] = (N154)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                          (N155)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                          (N156)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                          (N157)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                          (N158)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                          (N159)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                          (N160)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                          (N161)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                          (N162)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                          (N163)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                          (N164)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                          (N165)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                          (N166)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                          (N167)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                          (N168)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                          (N169)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                          (N170)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                          (N171)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                          (N172)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                          (N173)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                          (N174)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                          (N175)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                          (N176)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                          (N177)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                          (N178)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                          (N179)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                          (N180)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                          (N181)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                          (N182)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                          (N183)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                          (N184)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                          (N185)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                          (N186)? data_o[511:496] : 
                          (N187)? data_o[495:480] : 
                          (N188)? data_o[479:464] : 
                          (N189)? data_o[463:448] : 
                          (N190)? data_o[447:432] : 
                          (N191)? data_o[431:416] : 
                          (N192)? data_o[415:400] : 
                          (N193)? data_o[399:384] : 
                          (N194)? data_o[383:368] : 
                          (N195)? data_o[367:352] : 
                          (N196)? data_o[351:336] : 
                          (N197)? data_o[335:320] : 
                          (N198)? data_o[319:304] : 
                          (N199)? data_o[303:288] : 
                          (N200)? data_o[287:272] : 
                          (N201)? data_o[271:256] : 
                          (N202)? data_o[255:240] : 
                          (N203)? data_o[239:224] : 
                          (N204)? data_o[223:208] : 
                          (N205)? data_o[207:192] : 
                          (N206)? data_o[191:176] : 
                          (N207)? data_o[175:160] : 
                          (N208)? data_o[159:144] : 
                          (N209)? data_o[143:128] : 
                          (N210)? data_o[127:112] : 
                          (N211)? data_o[111:96] : 
                          (N212)? data_o[95:80] : 
                          (N213)? data_o[79:64] : 
                          (N214)? data_o[63:48] : 1'b0;
  assign data_nn[79:64] = (N155)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                          (N156)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                          (N157)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                          (N158)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                          (N159)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                          (N160)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                          (N161)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                          (N162)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                          (N163)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                          (N164)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                          (N165)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                          (N166)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                          (N167)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                          (N168)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                          (N169)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                          (N170)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                          (N171)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                          (N172)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                          (N173)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                          (N174)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                          (N175)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                          (N176)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                          (N177)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                          (N178)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                          (N179)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                          (N180)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                          (N181)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                          (N182)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                          (N183)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                          (N184)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                          (N185)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                          (N186)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                          (N187)? data_o[511:496] : 
                          (N188)? data_o[495:480] : 
                          (N189)? data_o[479:464] : 
                          (N190)? data_o[463:448] : 
                          (N191)? data_o[447:432] : 
                          (N192)? data_o[431:416] : 
                          (N193)? data_o[415:400] : 
                          (N194)? data_o[399:384] : 
                          (N195)? data_o[383:368] : 
                          (N196)? data_o[367:352] : 
                          (N197)? data_o[351:336] : 
                          (N198)? data_o[335:320] : 
                          (N199)? data_o[319:304] : 
                          (N200)? data_o[303:288] : 
                          (N201)? data_o[287:272] : 
                          (N202)? data_o[271:256] : 
                          (N203)? data_o[255:240] : 
                          (N204)? data_o[239:224] : 
                          (N205)? data_o[223:208] : 
                          (N206)? data_o[207:192] : 
                          (N207)? data_o[191:176] : 
                          (N208)? data_o[175:160] : 
                          (N209)? data_o[159:144] : 
                          (N210)? data_o[143:128] : 
                          (N211)? data_o[127:112] : 
                          (N212)? data_o[111:96] : 
                          (N213)? data_o[95:80] : 
                          (N214)? data_o[79:64] : 1'b0;
  assign data_nn[95:80] = (N156)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                          (N157)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                          (N158)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                          (N159)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                          (N160)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                          (N161)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                          (N162)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                          (N163)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                          (N164)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                          (N165)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                          (N166)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                          (N167)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                          (N168)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                          (N169)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                          (N170)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                          (N171)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                          (N172)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                          (N173)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                          (N174)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                          (N175)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                          (N176)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                          (N177)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                          (N178)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                          (N179)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                          (N180)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                          (N181)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                          (N182)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                          (N183)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                          (N184)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                          (N185)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                          (N186)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                          (N187)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                          (N188)? data_o[511:496] : 
                          (N189)? data_o[495:480] : 
                          (N190)? data_o[479:464] : 
                          (N191)? data_o[463:448] : 
                          (N192)? data_o[447:432] : 
                          (N193)? data_o[431:416] : 
                          (N194)? data_o[415:400] : 
                          (N195)? data_o[399:384] : 
                          (N196)? data_o[383:368] : 
                          (N197)? data_o[367:352] : 
                          (N198)? data_o[351:336] : 
                          (N199)? data_o[335:320] : 
                          (N200)? data_o[319:304] : 
                          (N201)? data_o[303:288] : 
                          (N202)? data_o[287:272] : 
                          (N203)? data_o[271:256] : 
                          (N204)? data_o[255:240] : 
                          (N205)? data_o[239:224] : 
                          (N206)? data_o[223:208] : 
                          (N207)? data_o[207:192] : 
                          (N208)? data_o[191:176] : 
                          (N209)? data_o[175:160] : 
                          (N210)? data_o[159:144] : 
                          (N211)? data_o[143:128] : 
                          (N212)? data_o[127:112] : 
                          (N213)? data_o[111:96] : 
                          (N214)? data_o[95:80] : 1'b0;
  assign data_nn[111:96] = (N157)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                           (N158)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                           (N159)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                           (N160)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                           (N161)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                           (N162)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                           (N163)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                           (N164)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                           (N165)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                           (N166)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                           (N167)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                           (N168)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                           (N169)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                           (N170)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                           (N171)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                           (N172)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                           (N173)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                           (N174)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                           (N175)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                           (N176)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                           (N177)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                           (N178)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                           (N179)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                           (N180)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                           (N181)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                           (N182)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                           (N183)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                           (N184)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                           (N185)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                           (N186)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                           (N187)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                           (N188)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                           (N189)? data_o[511:496] : 
                           (N190)? data_o[495:480] : 
                           (N191)? data_o[479:464] : 
                           (N192)? data_o[463:448] : 
                           (N193)? data_o[447:432] : 
                           (N194)? data_o[431:416] : 
                           (N195)? data_o[415:400] : 
                           (N196)? data_o[399:384] : 
                           (N197)? data_o[383:368] : 
                           (N198)? data_o[367:352] : 
                           (N199)? data_o[351:336] : 
                           (N200)? data_o[335:320] : 
                           (N201)? data_o[319:304] : 
                           (N202)? data_o[303:288] : 
                           (N203)? data_o[287:272] : 
                           (N204)? data_o[271:256] : 
                           (N205)? data_o[255:240] : 
                           (N206)? data_o[239:224] : 
                           (N207)? data_o[223:208] : 
                           (N208)? data_o[207:192] : 
                           (N209)? data_o[191:176] : 
                           (N210)? data_o[175:160] : 
                           (N211)? data_o[159:144] : 
                           (N212)? data_o[143:128] : 
                           (N213)? data_o[127:112] : 
                           (N214)? data_o[111:96] : 1'b0;
  assign data_nn[127:112] = (N215)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N159)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N160)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N161)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N162)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N216)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N217)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N218)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N219)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N167)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N168)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N169)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N170)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N220)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N221)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N222)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N223)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N175)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N176)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N177)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N178)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N224)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N225)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N226)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N227)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N228)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N229)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N230)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N231)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N232)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N233)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N234)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N235)? data_o[511:496] : 
                            (N236)? data_o[495:480] : 
                            (N237)? data_o[479:464] : 
                            (N238)? data_o[463:448] : 
                            (N239)? data_o[447:432] : 
                            (N240)? data_o[431:416] : 
                            (N241)? data_o[415:400] : 
                            (N242)? data_o[399:384] : 
                            (N243)? data_o[383:368] : 
                            (N244)? data_o[367:352] : 
                            (N245)? data_o[351:336] : 
                            (N246)? data_o[335:320] : 
                            (N247)? data_o[319:304] : 
                            (N248)? data_o[303:288] : 
                            (N249)? data_o[287:272] : 
                            (N250)? data_o[271:256] : 
                            (N251)? data_o[255:240] : 
                            (N252)? data_o[239:224] : 
                            (N253)? data_o[223:208] : 
                            (N254)? data_o[207:192] : 
                            (N255)? data_o[191:176] : 
                            (N256)? data_o[175:160] : 
                            (N257)? data_o[159:144] : 
                            (N258)? data_o[143:128] : 
                            (N259)? data_o[127:112] : 1'b0;
  assign N215 = N1346;
  assign N216 = N1351;
  assign N217 = N1352;
  assign N218 = N1353;
  assign N219 = N1354;
  assign N220 = N1359;
  assign N221 = N1360;
  assign N222 = N1361;
  assign N223 = N1362;
  assign N224 = N1367;
  assign N225 = N1368;
  assign N226 = N1369;
  assign N227 = N987;
  assign N228 = N986;
  assign N229 = N985;
  assign N230 = N984;
  assign N231 = N983;
  assign N232 = N982;
  assign N233 = N981;
  assign N234 = N980;
  assign N235 = N979;
  assign N236 = N978;
  assign N237 = N977;
  assign N238 = N976;
  assign N239 = N975;
  assign N240 = N974;
  assign N241 = N973;
  assign N242 = N972;
  assign N243 = N971;
  assign N244 = N970;
  assign N245 = N969;
  assign N246 = N968;
  assign N247 = N967;
  assign N248 = N966;
  assign N249 = N965;
  assign N250 = N964;
  assign N251 = N963;
  assign N252 = N962;
  assign N253 = N961;
  assign N254 = N960;
  assign N255 = N959;
  assign N256 = N958;
  assign N257 = N957;
  assign N258 = N956;
  assign N259 = N955;
  assign data_nn[143:128] = (N159)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N160)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N161)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N162)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N216)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N217)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N218)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N219)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N167)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N168)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N169)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N170)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N220)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N221)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N222)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N223)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N175)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N176)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N177)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N178)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N224)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N225)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N226)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N227)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N228)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N229)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N230)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N231)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N232)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N233)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N234)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N235)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N236)? data_o[511:496] : 
                            (N237)? data_o[495:480] : 
                            (N238)? data_o[479:464] : 
                            (N239)? data_o[463:448] : 
                            (N240)? data_o[447:432] : 
                            (N241)? data_o[431:416] : 
                            (N242)? data_o[415:400] : 
                            (N243)? data_o[399:384] : 
                            (N244)? data_o[383:368] : 
                            (N245)? data_o[367:352] : 
                            (N246)? data_o[351:336] : 
                            (N247)? data_o[335:320] : 
                            (N248)? data_o[319:304] : 
                            (N249)? data_o[303:288] : 
                            (N250)? data_o[287:272] : 
                            (N251)? data_o[271:256] : 
                            (N252)? data_o[255:240] : 
                            (N253)? data_o[239:224] : 
                            (N254)? data_o[223:208] : 
                            (N255)? data_o[207:192] : 
                            (N256)? data_o[191:176] : 
                            (N257)? data_o[175:160] : 
                            (N258)? data_o[159:144] : 
                            (N259)? data_o[143:128] : 1'b0;
  assign data_nn[159:144] = (N160)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N161)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N162)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N216)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N217)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N218)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N219)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N167)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N168)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N169)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N170)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N220)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N221)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N222)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N223)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N175)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N176)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N177)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N178)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N224)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N225)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N226)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N227)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N228)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N229)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N230)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N231)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N232)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N233)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N234)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N235)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N236)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N237)? data_o[511:496] : 
                            (N238)? data_o[495:480] : 
                            (N239)? data_o[479:464] : 
                            (N240)? data_o[463:448] : 
                            (N241)? data_o[447:432] : 
                            (N242)? data_o[431:416] : 
                            (N243)? data_o[415:400] : 
                            (N244)? data_o[399:384] : 
                            (N245)? data_o[383:368] : 
                            (N246)? data_o[367:352] : 
                            (N247)? data_o[351:336] : 
                            (N248)? data_o[335:320] : 
                            (N249)? data_o[319:304] : 
                            (N250)? data_o[303:288] : 
                            (N251)? data_o[287:272] : 
                            (N252)? data_o[271:256] : 
                            (N253)? data_o[255:240] : 
                            (N254)? data_o[239:224] : 
                            (N255)? data_o[223:208] : 
                            (N256)? data_o[207:192] : 
                            (N257)? data_o[191:176] : 
                            (N258)? data_o[175:160] : 
                            (N259)? data_o[159:144] : 1'b0;
  assign data_nn[175:160] = (N161)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N162)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N216)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N217)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N218)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N219)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N167)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N168)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N169)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N170)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N220)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N221)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N222)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N223)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N175)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N176)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N177)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N178)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N224)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N225)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N226)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N227)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N228)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N229)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N230)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N231)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N232)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N233)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N234)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N235)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N236)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N237)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N238)? data_o[511:496] : 
                            (N239)? data_o[495:480] : 
                            (N240)? data_o[479:464] : 
                            (N241)? data_o[463:448] : 
                            (N242)? data_o[447:432] : 
                            (N243)? data_o[431:416] : 
                            (N244)? data_o[415:400] : 
                            (N245)? data_o[399:384] : 
                            (N246)? data_o[383:368] : 
                            (N247)? data_o[367:352] : 
                            (N248)? data_o[351:336] : 
                            (N249)? data_o[335:320] : 
                            (N250)? data_o[319:304] : 
                            (N251)? data_o[303:288] : 
                            (N252)? data_o[287:272] : 
                            (N253)? data_o[271:256] : 
                            (N254)? data_o[255:240] : 
                            (N255)? data_o[239:224] : 
                            (N256)? data_o[223:208] : 
                            (N257)? data_o[207:192] : 
                            (N258)? data_o[191:176] : 
                            (N259)? data_o[175:160] : 1'b0;
  assign data_nn[191:176] = (N162)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N216)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N217)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N218)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N219)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N167)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N168)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N169)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N170)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N220)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N221)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N222)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N223)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N175)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N176)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N177)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N178)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N224)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N225)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N226)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N227)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N228)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N229)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N230)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N231)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N232)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N233)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N234)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N235)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N236)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N237)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N238)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N239)? data_o[511:496] : 
                            (N240)? data_o[495:480] : 
                            (N241)? data_o[479:464] : 
                            (N242)? data_o[463:448] : 
                            (N243)? data_o[447:432] : 
                            (N244)? data_o[431:416] : 
                            (N245)? data_o[415:400] : 
                            (N246)? data_o[399:384] : 
                            (N247)? data_o[383:368] : 
                            (N248)? data_o[367:352] : 
                            (N249)? data_o[351:336] : 
                            (N250)? data_o[335:320] : 
                            (N251)? data_o[319:304] : 
                            (N252)? data_o[303:288] : 
                            (N253)? data_o[287:272] : 
                            (N254)? data_o[271:256] : 
                            (N255)? data_o[255:240] : 
                            (N256)? data_o[239:224] : 
                            (N257)? data_o[223:208] : 
                            (N258)? data_o[207:192] : 
                            (N259)? data_o[191:176] : 1'b0;
  assign data_nn[207:192] = (N260)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N261)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N262)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N263)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N264)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N265)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N266)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N267)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N268)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N269)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N270)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N271)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N272)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N273)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N274)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N275)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N276)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N277)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N278)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N279)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N280)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N281)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N282)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N283)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N232)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N233)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N234)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N235)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N284)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N285)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N286)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N287)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N240)? data_o[511:496] : 
                            (N241)? data_o[495:480] : 
                            (N242)? data_o[479:464] : 
                            (N243)? data_o[463:448] : 
                            (N288)? data_o[447:432] : 
                            (N289)? data_o[431:416] : 
                            (N290)? data_o[415:400] : 
                            (N291)? data_o[399:384] : 
                            (N248)? data_o[383:368] : 
                            (N249)? data_o[367:352] : 
                            (N250)? data_o[351:336] : 
                            (N251)? data_o[335:320] : 
                            (N292)? data_o[319:304] : 
                            (N293)? data_o[303:288] : 
                            (N294)? data_o[287:272] : 
                            (N295)? data_o[271:256] : 
                            (N256)? data_o[255:240] : 
                            (N257)? data_o[239:224] : 
                            (N258)? data_o[223:208] : 
                            (N259)? data_o[207:192] : 1'b0;
  assign N260 = N1267;
  assign N261 = N1268;
  assign N262 = N1269;
  assign N263 = N1270;
  assign N264 = N1305;
  assign N265 = N1306;
  assign N266 = N1307;
  assign N267 = N1308;
  assign N268 = N865;
  assign N269 = N864;
  assign N270 = N863;
  assign N271 = N862;
  assign N272 = N1313;
  assign N273 = N1314;
  assign N274 = N1315;
  assign N275 = N1316;
  assign N276 = N861;
  assign N277 = N860;
  assign N278 = N859;
  assign N279 = N858;
  assign N280 = N857;
  assign N281 = N856;
  assign N282 = N855;
  assign N283 = N854;
  assign N284 = N853;
  assign N285 = N852;
  assign N286 = N851;
  assign N287 = N850;
  assign N288 = N849;
  assign N289 = N848;
  assign N290 = N847;
  assign N291 = N846;
  assign N292 = N845;
  assign N293 = N844;
  assign N294 = N843;
  assign N295 = N842;
  assign data_nn[223:208] = (N261)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N262)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N263)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N264)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N265)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N266)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N267)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N268)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N269)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N270)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N271)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N272)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N273)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N274)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N275)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N276)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N277)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N278)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N279)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N280)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N281)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N282)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N283)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N232)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N233)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N234)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N235)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N284)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N285)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N286)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N287)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N240)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N241)? data_o[511:496] : 
                            (N242)? data_o[495:480] : 
                            (N243)? data_o[479:464] : 
                            (N288)? data_o[463:448] : 
                            (N289)? data_o[447:432] : 
                            (N290)? data_o[431:416] : 
                            (N291)? data_o[415:400] : 
                            (N248)? data_o[399:384] : 
                            (N249)? data_o[383:368] : 
                            (N250)? data_o[367:352] : 
                            (N251)? data_o[351:336] : 
                            (N292)? data_o[335:320] : 
                            (N293)? data_o[319:304] : 
                            (N294)? data_o[303:288] : 
                            (N295)? data_o[287:272] : 
                            (N256)? data_o[271:256] : 
                            (N257)? data_o[255:240] : 
                            (N258)? data_o[239:224] : 
                            (N259)? data_o[223:208] : 1'b0;
  assign data_nn[239:224] = (N262)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N263)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N264)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N265)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N266)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N267)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N268)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N269)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N270)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N271)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N272)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N273)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N274)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N275)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N276)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N277)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N278)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N279)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N280)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N281)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N282)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N283)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N232)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N233)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N234)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N235)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N284)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N285)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N286)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N287)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N240)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N241)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N242)? data_o[511:496] : 
                            (N243)? data_o[495:480] : 
                            (N288)? data_o[479:464] : 
                            (N289)? data_o[463:448] : 
                            (N290)? data_o[447:432] : 
                            (N291)? data_o[431:416] : 
                            (N248)? data_o[415:400] : 
                            (N249)? data_o[399:384] : 
                            (N250)? data_o[383:368] : 
                            (N251)? data_o[367:352] : 
                            (N292)? data_o[351:336] : 
                            (N293)? data_o[335:320] : 
                            (N294)? data_o[319:304] : 
                            (N295)? data_o[303:288] : 
                            (N256)? data_o[287:272] : 
                            (N257)? data_o[271:256] : 
                            (N258)? data_o[255:240] : 
                            (N259)? data_o[239:224] : 1'b0;
  assign data_nn[255:240] = (N263)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N264)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N265)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N266)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N267)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N268)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N269)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N270)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N271)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N272)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N273)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N274)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N275)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N276)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N277)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N278)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N279)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N280)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N281)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N282)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N283)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N232)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N233)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N234)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N235)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N284)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N285)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N286)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N287)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N240)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N241)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N242)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N243)? data_o[511:496] : 
                            (N288)? data_o[495:480] : 
                            (N289)? data_o[479:464] : 
                            (N290)? data_o[463:448] : 
                            (N291)? data_o[447:432] : 
                            (N248)? data_o[431:416] : 
                            (N249)? data_o[415:400] : 
                            (N250)? data_o[399:384] : 
                            (N251)? data_o[383:368] : 
                            (N292)? data_o[367:352] : 
                            (N293)? data_o[351:336] : 
                            (N294)? data_o[335:320] : 
                            (N295)? data_o[319:304] : 
                            (N256)? data_o[303:288] : 
                            (N257)? data_o[287:272] : 
                            (N258)? data_o[271:256] : 
                            (N259)? data_o[255:240] : 1'b0;
  assign data_nn[271:256] = (N264)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N265)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N266)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N267)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N268)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N269)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N270)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N271)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N272)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N273)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N274)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N275)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N276)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N277)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N278)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N279)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N280)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N281)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N282)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N283)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N232)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N233)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N234)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N235)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N284)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N285)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N286)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N287)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N240)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N241)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N242)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N243)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N288)? data_o[511:496] : 
                            (N289)? data_o[495:480] : 
                            (N290)? data_o[479:464] : 
                            (N291)? data_o[463:448] : 
                            (N248)? data_o[447:432] : 
                            (N249)? data_o[431:416] : 
                            (N250)? data_o[415:400] : 
                            (N251)? data_o[399:384] : 
                            (N292)? data_o[383:368] : 
                            (N293)? data_o[367:352] : 
                            (N294)? data_o[351:336] : 
                            (N295)? data_o[335:320] : 
                            (N256)? data_o[319:304] : 
                            (N257)? data_o[303:288] : 
                            (N258)? data_o[287:272] : 
                            (N259)? data_o[271:256] : 1'b0;
  assign data_nn[287:272] = (N265)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N266)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N267)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N268)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N269)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N270)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N271)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N272)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N273)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N274)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N275)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N276)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N277)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N278)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N279)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N280)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N281)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N282)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N283)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N232)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N233)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N234)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N235)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N284)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N285)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N286)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N287)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N240)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N241)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N242)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N243)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N288)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N289)? data_o[511:496] : 
                            (N290)? data_o[495:480] : 
                            (N291)? data_o[479:464] : 
                            (N248)? data_o[463:448] : 
                            (N249)? data_o[447:432] : 
                            (N250)? data_o[431:416] : 
                            (N251)? data_o[415:400] : 
                            (N292)? data_o[399:384] : 
                            (N293)? data_o[383:368] : 
                            (N294)? data_o[367:352] : 
                            (N295)? data_o[351:336] : 
                            (N256)? data_o[335:320] : 
                            (N257)? data_o[319:304] : 
                            (N258)? data_o[303:288] : 
                            (N259)? data_o[287:272] : 1'b0;
  assign data_nn[303:288] = (N266)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N267)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N296)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N297)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N298)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N299)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N272)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N273)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N274)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N275)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N300)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N301)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N302)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N303)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N304)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N305)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N306)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N307)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N308)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N309)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N310)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N311)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N312)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N313)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N314)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N315)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N316)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N317)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N318)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N319)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N320)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N321)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N322)? data_o[511:496] : 
                            (N323)? data_o[495:480] : 
                            (N324)? data_o[479:464] : 
                            (N325)? data_o[463:448] : 
                            (N326)? data_o[447:432] : 
                            (N327)? data_o[431:416] : 
                            (N328)? data_o[415:400] : 
                            (N329)? data_o[399:384] : 
                            (N330)? data_o[383:368] : 
                            (N331)? data_o[367:352] : 
                            (N332)? data_o[351:336] : 
                            (N333)? data_o[335:320] : 
                            (N334)? data_o[319:304] : 
                            (N335)? data_o[303:288] : 1'b0;
  assign N296 = N1309;
  assign N297 = N1310;
  assign N298 = N1311;
  assign N299 = N1312;
  assign N300 = N1317;
  assign N301 = N1318;
  assign N302 = N954;
  assign N303 = N953;
  assign N304 = N952;
  assign N305 = N951;
  assign N306 = N950;
  assign N307 = N949;
  assign N308 = N948;
  assign N309 = N947;
  assign N310 = N946;
  assign N311 = N945;
  assign N312 = N944;
  assign N313 = N943;
  assign N314 = N942;
  assign N315 = N941;
  assign N316 = N940;
  assign N317 = N939;
  assign N318 = N938;
  assign N319 = N937;
  assign N320 = N936;
  assign N321 = N935;
  assign N322 = N934;
  assign N323 = N933;
  assign N324 = N932;
  assign N325 = N931;
  assign N326 = N930;
  assign N327 = N929;
  assign N328 = N928;
  assign N329 = N927;
  assign N330 = N926;
  assign N331 = N925;
  assign N332 = N924;
  assign N333 = N923;
  assign N334 = N922;
  assign N335 = N921;
  assign data_nn[319:304] = (N267)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N296)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N297)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N298)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N299)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N272)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N273)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N274)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N275)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N300)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N301)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N302)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N303)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N304)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N305)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N306)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N307)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N308)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N309)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N310)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N311)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N312)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N313)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N314)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N315)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N316)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N317)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N318)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N319)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N320)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N321)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N322)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N323)? data_o[511:496] : 
                            (N324)? data_o[495:480] : 
                            (N325)? data_o[479:464] : 
                            (N326)? data_o[463:448] : 
                            (N327)? data_o[447:432] : 
                            (N328)? data_o[431:416] : 
                            (N329)? data_o[415:400] : 
                            (N330)? data_o[399:384] : 
                            (N331)? data_o[383:368] : 
                            (N332)? data_o[367:352] : 
                            (N333)? data_o[351:336] : 
                            (N334)? data_o[335:320] : 
                            (N335)? data_o[319:304] : 1'b0;
  assign data_nn[335:320] = (N296)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N297)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N298)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N299)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N272)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N273)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N274)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N275)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N300)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N301)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N302)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N303)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N304)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N305)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N306)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N307)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N308)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N309)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N310)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N311)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N312)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N313)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N314)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N315)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N316)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N317)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N318)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N319)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N320)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N321)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N322)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N323)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N324)? data_o[511:496] : 
                            (N325)? data_o[495:480] : 
                            (N326)? data_o[479:464] : 
                            (N327)? data_o[463:448] : 
                            (N328)? data_o[447:432] : 
                            (N329)? data_o[431:416] : 
                            (N330)? data_o[415:400] : 
                            (N331)? data_o[399:384] : 
                            (N332)? data_o[383:368] : 
                            (N333)? data_o[367:352] : 
                            (N334)? data_o[351:336] : 
                            (N335)? data_o[335:320] : 1'b0;
  assign data_nn[351:336] = (N297)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N298)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N299)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N272)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N273)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N274)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N275)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N300)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N301)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N302)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N303)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N304)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N305)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N306)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N307)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N308)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N309)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N310)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N311)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N312)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N313)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N314)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N315)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N316)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N317)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N318)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N319)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N320)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N321)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N322)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N323)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N324)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N325)? data_o[511:496] : 
                            (N326)? data_o[495:480] : 
                            (N327)? data_o[479:464] : 
                            (N328)? data_o[463:448] : 
                            (N329)? data_o[447:432] : 
                            (N330)? data_o[431:416] : 
                            (N331)? data_o[415:400] : 
                            (N332)? data_o[399:384] : 
                            (N333)? data_o[383:368] : 
                            (N334)? data_o[367:352] : 
                            (N335)? data_o[351:336] : 1'b0;
  assign data_nn[367:352] = (N298)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N299)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N272)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N273)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N274)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N275)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N300)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N301)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N302)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N303)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N304)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N305)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N306)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N307)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N308)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N309)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N310)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N311)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N312)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N313)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N314)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N315)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N316)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N317)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N318)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N319)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N320)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N321)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N322)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N323)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N324)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N325)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N326)? data_o[511:496] : 
                            (N327)? data_o[495:480] : 
                            (N328)? data_o[479:464] : 
                            (N329)? data_o[463:448] : 
                            (N330)? data_o[447:432] : 
                            (N331)? data_o[431:416] : 
                            (N332)? data_o[415:400] : 
                            (N333)? data_o[399:384] : 
                            (N334)? data_o[383:368] : 
                            (N335)? data_o[367:352] : 1'b0;
  assign data_nn[383:368] = (N336)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N337)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N338)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N339)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N340)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N341)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N342)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N343)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N344)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N345)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N346)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N347)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N348)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N308)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N309)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N310)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N311)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N349)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N350)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N351)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N352)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N316)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N317)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N318)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N319)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N353)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N354)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N355)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N356)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N324)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N325)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N326)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N327)? data_o[511:496] : 
                            (N357)? data_o[495:480] : 
                            (N358)? data_o[479:464] : 
                            (N359)? data_o[463:448] : 
                            (N360)? data_o[447:432] : 
                            (N332)? data_o[431:416] : 
                            (N333)? data_o[415:400] : 
                            (N334)? data_o[399:384] : 
                            (N335)? data_o[383:368] : 1'b0;
  assign N336 = N1271;
  assign N337 = N1286;
  assign N338 = N1287;
  assign N339 = N1288;
  assign N340 = N1289;
  assign N341 = N885;
  assign N342 = N884;
  assign N343 = N883;
  assign N344 = N882;
  assign N345 = N881;
  assign N346 = N880;
  assign N347 = N879;
  assign N348 = N878;
  assign N349 = N877;
  assign N350 = N876;
  assign N351 = N875;
  assign N352 = N874;
  assign N353 = N873;
  assign N354 = N872;
  assign N355 = N871;
  assign N356 = N870;
  assign N357 = N869;
  assign N358 = N868;
  assign N359 = N867;
  assign N360 = N866;
  assign data_nn[399:384] = (N337)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N338)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N339)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N340)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N341)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N342)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N343)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N344)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N345)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N346)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N347)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N348)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N308)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N309)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N310)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N311)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N349)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N350)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N351)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N352)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N316)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N317)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N318)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N319)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N353)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N354)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N355)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N356)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N324)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N325)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N326)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N327)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N357)? data_o[511:496] : 
                            (N358)? data_o[495:480] : 
                            (N359)? data_o[479:464] : 
                            (N360)? data_o[463:448] : 
                            (N332)? data_o[447:432] : 
                            (N333)? data_o[431:416] : 
                            (N334)? data_o[415:400] : 
                            (N335)? data_o[399:384] : 1'b0;
  assign data_nn[415:400] = (N338)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N339)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N340)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N341)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N342)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N343)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N344)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N345)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N346)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N347)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N348)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N308)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N309)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N310)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N311)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N349)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N350)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N351)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N352)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N316)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N317)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N318)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N319)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N353)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N354)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N355)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N356)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N324)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N325)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N326)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N327)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N357)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N358)? data_o[511:496] : 
                            (N359)? data_o[495:480] : 
                            (N360)? data_o[479:464] : 
                            (N332)? data_o[463:448] : 
                            (N333)? data_o[447:432] : 
                            (N334)? data_o[431:416] : 
                            (N335)? data_o[415:400] : 1'b0;
  assign data_nn[431:416] = (N339)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N340)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N341)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N342)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N343)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N344)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N345)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N346)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N347)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N348)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N308)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N309)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N310)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N311)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N349)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N350)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N351)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N352)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N316)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N317)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N318)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N319)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N353)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N354)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N355)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N356)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N324)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N325)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N326)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N327)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N357)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N358)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N359)? data_o[511:496] : 
                            (N360)? data_o[495:480] : 
                            (N332)? data_o[479:464] : 
                            (N333)? data_o[463:448] : 
                            (N334)? data_o[447:432] : 
                            (N335)? data_o[431:416] : 1'b0;
  assign data_nn[447:432] = (N340)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N341)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N342)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N343)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N344)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N345)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N346)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N347)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N348)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N308)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N309)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N310)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N311)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N349)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N350)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N351)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N352)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N316)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N317)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N318)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N319)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N353)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N354)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N355)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N356)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N324)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N325)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N326)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N327)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N357)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N358)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N359)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N360)? data_o[511:496] : 
                            (N332)? data_o[495:480] : 
                            (N333)? data_o[479:464] : 
                            (N334)? data_o[463:448] : 
                            (N335)? data_o[447:432] : 1'b0;
  assign data_nn[463:448] = (N341)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N342)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N343)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N344)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N345)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N346)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N347)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N348)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N308)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N309)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N310)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N311)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N349)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N350)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N351)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N352)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N316)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N317)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N318)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N319)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N353)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N354)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N355)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N356)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N324)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N325)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N326)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N327)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N357)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N358)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N359)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N360)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N332)? data_o[511:496] : 
                            (N333)? data_o[495:480] : 
                            (N334)? data_o[479:464] : 
                            (N335)? data_o[463:448] : 1'b0;
  assign data_nn[479:464] = (N361)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N362)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N363)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N364)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N365)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N366)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N367)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N368)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N369)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N370)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N371)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N372)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N373)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N374)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N375)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N376)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N377)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N378)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N379)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N380)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N381)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N382)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N383)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N384)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N385)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N386)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N387)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N388)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N389)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N390)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N391)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N392)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N393)? data_o[511:496] : 
                            (N394)? data_o[495:480] : 
                            (N395)? data_o[479:464] : 1'b0;
  assign N361 = N920;
  assign N362 = N919;
  assign N363 = N918;
  assign N364 = N917;
  assign N365 = N916;
  assign N366 = N915;
  assign N367 = N914;
  assign N368 = N913;
  assign N369 = N912;
  assign N370 = N911;
  assign N371 = N910;
  assign N372 = N909;
  assign N373 = N908;
  assign N374 = N907;
  assign N375 = N906;
  assign N376 = N905;
  assign N377 = N904;
  assign N378 = N903;
  assign N379 = N902;
  assign N380 = N901;
  assign N381 = N900;
  assign N382 = N899;
  assign N383 = N898;
  assign N384 = N897;
  assign N385 = N896;
  assign N386 = N895;
  assign N387 = N894;
  assign N388 = N893;
  assign N389 = N892;
  assign N390 = N891;
  assign N391 = N890;
  assign N392 = N889;
  assign N393 = N888;
  assign N394 = N887;
  assign N395 = N886;
  assign data_nn[495:480] = (N302)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N303)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N304)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N305)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N306)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N307)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N308)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N309)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N310)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N311)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N312)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N313)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N314)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N315)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N316)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N317)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N318)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N319)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N320)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N321)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N322)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N323)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N324)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N325)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N326)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N327)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N328)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N329)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N330)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N331)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N332)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N333)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N334)? data_o[511:496] : 
                            (N335)? data_o[495:480] : 1'b0;
  assign data_nn[511:496] = (N227)? { data_n_63__15_, data_n_63__14_, data_n_63__13_, data_n_63__12_, data_n_63__11_, data_n_63__10_, data_n_63__9_, data_n_63__8_, data_n_63__7_, data_n_63__6_, data_n_63__5_, data_n_63__4_, data_n_63__3_, data_n_63__2_, data_n_63__1_, data_n_63__0_ } : 
                            (N228)? { data_n_62__15_, data_n_62__14_, data_n_62__13_, data_n_62__12_, data_n_62__11_, data_n_62__10_, data_n_62__9_, data_n_62__8_, data_n_62__7_, data_n_62__6_, data_n_62__5_, data_n_62__4_, data_n_62__3_, data_n_62__2_, data_n_62__1_, data_n_62__0_ } : 
                            (N229)? { data_n_61__15_, data_n_61__14_, data_n_61__13_, data_n_61__12_, data_n_61__11_, data_n_61__10_, data_n_61__9_, data_n_61__8_, data_n_61__7_, data_n_61__6_, data_n_61__5_, data_n_61__4_, data_n_61__3_, data_n_61__2_, data_n_61__1_, data_n_61__0_ } : 
                            (N230)? { data_n_60__15_, data_n_60__14_, data_n_60__13_, data_n_60__12_, data_n_60__11_, data_n_60__10_, data_n_60__9_, data_n_60__8_, data_n_60__7_, data_n_60__6_, data_n_60__5_, data_n_60__4_, data_n_60__3_, data_n_60__2_, data_n_60__1_, data_n_60__0_ } : 
                            (N231)? { data_n_59__15_, data_n_59__14_, data_n_59__13_, data_n_59__12_, data_n_59__11_, data_n_59__10_, data_n_59__9_, data_n_59__8_, data_n_59__7_, data_n_59__6_, data_n_59__5_, data_n_59__4_, data_n_59__3_, data_n_59__2_, data_n_59__1_, data_n_59__0_ } : 
                            (N232)? { data_n_58__15_, data_n_58__14_, data_n_58__13_, data_n_58__12_, data_n_58__11_, data_n_58__10_, data_n_58__9_, data_n_58__8_, data_n_58__7_, data_n_58__6_, data_n_58__5_, data_n_58__4_, data_n_58__3_, data_n_58__2_, data_n_58__1_, data_n_58__0_ } : 
                            (N233)? { data_n_57__15_, data_n_57__14_, data_n_57__13_, data_n_57__12_, data_n_57__11_, data_n_57__10_, data_n_57__9_, data_n_57__8_, data_n_57__7_, data_n_57__6_, data_n_57__5_, data_n_57__4_, data_n_57__3_, data_n_57__2_, data_n_57__1_, data_n_57__0_ } : 
                            (N234)? { data_n_56__15_, data_n_56__14_, data_n_56__13_, data_n_56__12_, data_n_56__11_, data_n_56__10_, data_n_56__9_, data_n_56__8_, data_n_56__7_, data_n_56__6_, data_n_56__5_, data_n_56__4_, data_n_56__3_, data_n_56__2_, data_n_56__1_, data_n_56__0_ } : 
                            (N235)? { data_n_55__15_, data_n_55__14_, data_n_55__13_, data_n_55__12_, data_n_55__11_, data_n_55__10_, data_n_55__9_, data_n_55__8_, data_n_55__7_, data_n_55__6_, data_n_55__5_, data_n_55__4_, data_n_55__3_, data_n_55__2_, data_n_55__1_, data_n_55__0_ } : 
                            (N236)? { data_n_54__15_, data_n_54__14_, data_n_54__13_, data_n_54__12_, data_n_54__11_, data_n_54__10_, data_n_54__9_, data_n_54__8_, data_n_54__7_, data_n_54__6_, data_n_54__5_, data_n_54__4_, data_n_54__3_, data_n_54__2_, data_n_54__1_, data_n_54__0_ } : 
                            (N237)? { data_n_53__15_, data_n_53__14_, data_n_53__13_, data_n_53__12_, data_n_53__11_, data_n_53__10_, data_n_53__9_, data_n_53__8_, data_n_53__7_, data_n_53__6_, data_n_53__5_, data_n_53__4_, data_n_53__3_, data_n_53__2_, data_n_53__1_, data_n_53__0_ } : 
                            (N238)? { data_n_52__15_, data_n_52__14_, data_n_52__13_, data_n_52__12_, data_n_52__11_, data_n_52__10_, data_n_52__9_, data_n_52__8_, data_n_52__7_, data_n_52__6_, data_n_52__5_, data_n_52__4_, data_n_52__3_, data_n_52__2_, data_n_52__1_, data_n_52__0_ } : 
                            (N239)? { data_n_51__15_, data_n_51__14_, data_n_51__13_, data_n_51__12_, data_n_51__11_, data_n_51__10_, data_n_51__9_, data_n_51__8_, data_n_51__7_, data_n_51__6_, data_n_51__5_, data_n_51__4_, data_n_51__3_, data_n_51__2_, data_n_51__1_, data_n_51__0_ } : 
                            (N240)? { data_n_50__15_, data_n_50__14_, data_n_50__13_, data_n_50__12_, data_n_50__11_, data_n_50__10_, data_n_50__9_, data_n_50__8_, data_n_50__7_, data_n_50__6_, data_n_50__5_, data_n_50__4_, data_n_50__3_, data_n_50__2_, data_n_50__1_, data_n_50__0_ } : 
                            (N241)? { data_n_49__15_, data_n_49__14_, data_n_49__13_, data_n_49__12_, data_n_49__11_, data_n_49__10_, data_n_49__9_, data_n_49__8_, data_n_49__7_, data_n_49__6_, data_n_49__5_, data_n_49__4_, data_n_49__3_, data_n_49__2_, data_n_49__1_, data_n_49__0_ } : 
                            (N242)? { data_n_48__15_, data_n_48__14_, data_n_48__13_, data_n_48__12_, data_n_48__11_, data_n_48__10_, data_n_48__9_, data_n_48__8_, data_n_48__7_, data_n_48__6_, data_n_48__5_, data_n_48__4_, data_n_48__3_, data_n_48__2_, data_n_48__1_, data_n_48__0_ } : 
                            (N243)? { data_n_47__15_, data_n_47__14_, data_n_47__13_, data_n_47__12_, data_n_47__11_, data_n_47__10_, data_n_47__9_, data_n_47__8_, data_n_47__7_, data_n_47__6_, data_n_47__5_, data_n_47__4_, data_n_47__3_, data_n_47__2_, data_n_47__1_, data_n_47__0_ } : 
                            (N244)? { data_n_46__15_, data_n_46__14_, data_n_46__13_, data_n_46__12_, data_n_46__11_, data_n_46__10_, data_n_46__9_, data_n_46__8_, data_n_46__7_, data_n_46__6_, data_n_46__5_, data_n_46__4_, data_n_46__3_, data_n_46__2_, data_n_46__1_, data_n_46__0_ } : 
                            (N245)? { data_n_45__15_, data_n_45__14_, data_n_45__13_, data_n_45__12_, data_n_45__11_, data_n_45__10_, data_n_45__9_, data_n_45__8_, data_n_45__7_, data_n_45__6_, data_n_45__5_, data_n_45__4_, data_n_45__3_, data_n_45__2_, data_n_45__1_, data_n_45__0_ } : 
                            (N246)? { data_n_44__15_, data_n_44__14_, data_n_44__13_, data_n_44__12_, data_n_44__11_, data_n_44__10_, data_n_44__9_, data_n_44__8_, data_n_44__7_, data_n_44__6_, data_n_44__5_, data_n_44__4_, data_n_44__3_, data_n_44__2_, data_n_44__1_, data_n_44__0_ } : 
                            (N247)? { data_n_43__15_, data_n_43__14_, data_n_43__13_, data_n_43__12_, data_n_43__11_, data_n_43__10_, data_n_43__9_, data_n_43__8_, data_n_43__7_, data_n_43__6_, data_n_43__5_, data_n_43__4_, data_n_43__3_, data_n_43__2_, data_n_43__1_, data_n_43__0_ } : 
                            (N248)? { data_n_42__15_, data_n_42__14_, data_n_42__13_, data_n_42__12_, data_n_42__11_, data_n_42__10_, data_n_42__9_, data_n_42__8_, data_n_42__7_, data_n_42__6_, data_n_42__5_, data_n_42__4_, data_n_42__3_, data_n_42__2_, data_n_42__1_, data_n_42__0_ } : 
                            (N249)? { data_n_41__15_, data_n_41__14_, data_n_41__13_, data_n_41__12_, data_n_41__11_, data_n_41__10_, data_n_41__9_, data_n_41__8_, data_n_41__7_, data_n_41__6_, data_n_41__5_, data_n_41__4_, data_n_41__3_, data_n_41__2_, data_n_41__1_, data_n_41__0_ } : 
                            (N250)? { data_n_40__15_, data_n_40__14_, data_n_40__13_, data_n_40__12_, data_n_40__11_, data_n_40__10_, data_n_40__9_, data_n_40__8_, data_n_40__7_, data_n_40__6_, data_n_40__5_, data_n_40__4_, data_n_40__3_, data_n_40__2_, data_n_40__1_, data_n_40__0_ } : 
                            (N251)? { data_n_39__15_, data_n_39__14_, data_n_39__13_, data_n_39__12_, data_n_39__11_, data_n_39__10_, data_n_39__9_, data_n_39__8_, data_n_39__7_, data_n_39__6_, data_n_39__5_, data_n_39__4_, data_n_39__3_, data_n_39__2_, data_n_39__1_, data_n_39__0_ } : 
                            (N252)? { data_n_38__15_, data_n_38__14_, data_n_38__13_, data_n_38__12_, data_n_38__11_, data_n_38__10_, data_n_38__9_, data_n_38__8_, data_n_38__7_, data_n_38__6_, data_n_38__5_, data_n_38__4_, data_n_38__3_, data_n_38__2_, data_n_38__1_, data_n_38__0_ } : 
                            (N253)? { data_n_37__15_, data_n_37__14_, data_n_37__13_, data_n_37__12_, data_n_37__11_, data_n_37__10_, data_n_37__9_, data_n_37__8_, data_n_37__7_, data_n_37__6_, data_n_37__5_, data_n_37__4_, data_n_37__3_, data_n_37__2_, data_n_37__1_, data_n_37__0_ } : 
                            (N254)? { data_n_36__15_, data_n_36__14_, data_n_36__13_, data_n_36__12_, data_n_36__11_, data_n_36__10_, data_n_36__9_, data_n_36__8_, data_n_36__7_, data_n_36__6_, data_n_36__5_, data_n_36__4_, data_n_36__3_, data_n_36__2_, data_n_36__1_, data_n_36__0_ } : 
                            (N255)? { data_n_35__15_, data_n_35__14_, data_n_35__13_, data_n_35__12_, data_n_35__11_, data_n_35__10_, data_n_35__9_, data_n_35__8_, data_n_35__7_, data_n_35__6_, data_n_35__5_, data_n_35__4_, data_n_35__3_, data_n_35__2_, data_n_35__1_, data_n_35__0_ } : 
                            (N256)? { data_n_34__15_, data_n_34__14_, data_n_34__13_, data_n_34__12_, data_n_34__11_, data_n_34__10_, data_n_34__9_, data_n_34__8_, data_n_34__7_, data_n_34__6_, data_n_34__5_, data_n_34__4_, data_n_34__3_, data_n_34__2_, data_n_34__1_, data_n_34__0_ } : 
                            (N257)? { data_n_33__15_, data_n_33__14_, data_n_33__13_, data_n_33__12_, data_n_33__11_, data_n_33__10_, data_n_33__9_, data_n_33__8_, data_n_33__7_, data_n_33__6_, data_n_33__5_, data_n_33__4_, data_n_33__3_, data_n_33__2_, data_n_33__1_, data_n_33__0_ } : 
                            (N258)? { data_n_32__15_, data_n_32__14_, data_n_32__13_, data_n_32__12_, data_n_32__11_, data_n_32__10_, data_n_32__9_, data_n_32__8_, data_n_32__7_, data_n_32__6_, data_n_32__5_, data_n_32__4_, data_n_32__3_, data_n_32__2_, data_n_32__1_, data_n_32__0_ } : 
                            (N259)? data_o[511:496] : 1'b0;
  assign { N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988 } = (N396)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, valid_n } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                           (N731)? { valid_n[62:32], valid_o } : 1'b0;
  assign N396 = yumi_cnt_i[5];
  assign { N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051 } = (N397)? { N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004 } : 
                                                                                                                                                                                                                                                                                                                                                       (N698)? { N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988 } : 1'b0;
  assign N397 = yumi_cnt_i[4];
  assign { N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098 } = (N398)? { N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059 } : 
                                                                                                                                                                                                                                                                                               (N681)? { N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051 } : 1'b0;
  assign N398 = yumi_cnt_i[3];
  assign { N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137 } = (N399)? { N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102 } : 
                                                                                                                                                                                                                                                                   (N672)? { N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098 } : 1'b0;
  assign N399 = yumi_cnt_i[2];
  assign { N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172 } = (N400)? { N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139 } : 
                                                                                                                                                                                                                                                     (N667)? { N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137 } : 1'b0;
  assign N400 = yumi_cnt_i[1];
  assign valid_nn = (N401)? { N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173 } : 
                    (N666)? { N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172 } : 1'b0;
  assign N401 = yumi_cnt_i[0];
  assign ready_o = ~valid_r[31];
  assign N402 = valid_i & ready_o;
  assign N473 = ~N409;
  assign N474 = ~N410;
  assign N475 = ~N411;
  assign N476 = ~N412;
  assign N477 = ~N413;
  assign N478 = ~N414;
  assign N479 = ~N415;
  assign N480 = ~N416;
  assign N481 = ~N417;
  assign N482 = ~N418;
  assign N483 = ~N419;
  assign N484 = ~N420;
  assign N485 = ~N421;
  assign N486 = ~N422;
  assign N487 = ~N423;
  assign N488 = ~N424;
  assign N489 = ~N425;
  assign N490 = ~N426;
  assign N491 = ~N427;
  assign N492 = ~N428;
  assign N493 = ~N429;
  assign N494 = ~N430;
  assign N495 = ~N431;
  assign N496 = ~N432;
  assign N497 = ~N433;
  assign N498 = ~N434;
  assign N499 = ~N435;
  assign N500 = ~N436;
  assign N501 = ~N437;
  assign N502 = ~N438;
  assign N503 = ~N439;
  assign N504 = ~N440;
  assign N505 = ~N441;
  assign N506 = ~N442;
  assign N507 = ~N443;
  assign N508 = ~N444;
  assign N509 = ~N445;
  assign N510 = ~N446;
  assign N511 = ~N447;
  assign N512 = ~N448;
  assign N513 = ~N449;
  assign N514 = ~N450;
  assign N515 = ~N451;
  assign N516 = ~N452;
  assign N517 = ~N453;
  assign N518 = ~N454;
  assign N519 = ~N455;
  assign N520 = ~N456;
  assign N521 = ~N457;
  assign N522 = ~N458;
  assign N523 = ~N459;
  assign N524 = ~N460;
  assign N525 = ~N461;
  assign N526 = ~N462;
  assign N527 = ~N463;
  assign N528 = ~N464;
  assign N529 = ~N465;
  assign N530 = ~N466;
  assign N531 = ~N467;
  assign N532 = ~N468;
  assign N533 = ~N469;
  assign N534 = ~N470;
  assign N535 = ~N471;
  assign N536 = ~N472;
  assign N601 = valid_i & ready_o;
  assign N602 = ~N537;
  assign N603 = ~N538;
  assign N604 = ~N539;
  assign N605 = ~N540;
  assign N606 = ~N541;
  assign N607 = ~N542;
  assign N608 = ~N543;
  assign N609 = ~N544;
  assign N610 = ~N545;
  assign N611 = ~N546;
  assign N612 = ~N547;
  assign N613 = ~N548;
  assign N614 = ~N549;
  assign N615 = ~N550;
  assign N616 = ~N551;
  assign N617 = ~N552;
  assign N618 = ~N553;
  assign N619 = ~N554;
  assign N620 = ~N555;
  assign N621 = ~N556;
  assign N622 = ~N557;
  assign N623 = ~N558;
  assign N624 = ~N559;
  assign N625 = ~N560;
  assign N626 = ~N561;
  assign N627 = ~N562;
  assign N628 = ~N563;
  assign N629 = ~N564;
  assign N630 = ~N565;
  assign N631 = ~N566;
  assign N632 = ~N567;
  assign N633 = ~N568;
  assign N634 = ~N569;
  assign N635 = ~N570;
  assign N636 = ~N571;
  assign N637 = ~N572;
  assign N638 = ~N573;
  assign N639 = ~N574;
  assign N640 = ~N575;
  assign N641 = ~N576;
  assign N642 = ~N577;
  assign N643 = ~N578;
  assign N644 = ~N579;
  assign N645 = ~N580;
  assign N646 = ~N581;
  assign N647 = ~N582;
  assign N648 = ~N583;
  assign N649 = ~N584;
  assign N650 = ~N585;
  assign N651 = ~N586;
  assign N652 = ~N587;
  assign N653 = ~N588;
  assign N654 = ~N589;
  assign N655 = ~N590;
  assign N656 = ~N591;
  assign N657 = ~N592;
  assign N658 = ~N593;
  assign N659 = ~N594;
  assign N660 = ~N595;
  assign N661 = ~N596;
  assign N662 = ~N597;
  assign N663 = ~N598;
  assign N664 = ~N599;
  assign N665 = ~N600;
  assign N666 = ~yumi_cnt_i[0];
  assign N667 = ~yumi_cnt_i[1];
  assign N668 = N666 & N667;
  assign N669 = N666 & yumi_cnt_i[1];
  assign N670 = yumi_cnt_i[0] & N667;
  assign N671 = yumi_cnt_i[0] & yumi_cnt_i[1];
  assign N672 = ~yumi_cnt_i[2];
  assign N673 = N668 & N672;
  assign N674 = N668 & yumi_cnt_i[2];
  assign N675 = N670 & N672;
  assign N676 = N670 & yumi_cnt_i[2];
  assign N677 = N669 & N672;
  assign N678 = N669 & yumi_cnt_i[2];
  assign N679 = N671 & N672;
  assign N680 = N671 & yumi_cnt_i[2];
  assign N681 = ~yumi_cnt_i[3];
  assign N682 = N673 & N681;
  assign N683 = N673 & yumi_cnt_i[3];
  assign N684 = N675 & N681;
  assign N685 = N675 & yumi_cnt_i[3];
  assign N686 = N677 & N681;
  assign N687 = N677 & yumi_cnt_i[3];
  assign N688 = N679 & N681;
  assign N689 = N679 & yumi_cnt_i[3];
  assign N690 = N674 & N681;
  assign N691 = N674 & yumi_cnt_i[3];
  assign N692 = N676 & N681;
  assign N693 = N676 & yumi_cnt_i[3];
  assign N694 = N678 & N681;
  assign N695 = N678 & yumi_cnt_i[3];
  assign N696 = N680 & N681;
  assign N697 = N680 & yumi_cnt_i[3];
  assign N698 = ~yumi_cnt_i[4];
  assign N699 = N682 & N698;
  assign N700 = N682 & yumi_cnt_i[4];
  assign N701 = N684 & N698;
  assign N702 = N684 & yumi_cnt_i[4];
  assign N703 = N686 & N698;
  assign N704 = N686 & yumi_cnt_i[4];
  assign N705 = N688 & N698;
  assign N706 = N688 & yumi_cnt_i[4];
  assign N707 = N690 & N698;
  assign N708 = N690 & yumi_cnt_i[4];
  assign N709 = N692 & N698;
  assign N710 = N692 & yumi_cnt_i[4];
  assign N711 = N694 & N698;
  assign N712 = N694 & yumi_cnt_i[4];
  assign N713 = N696 & N698;
  assign N714 = N696 & yumi_cnt_i[4];
  assign N715 = N683 & N698;
  assign N716 = N683 & yumi_cnt_i[4];
  assign N717 = N685 & N698;
  assign N718 = N685 & yumi_cnt_i[4];
  assign N719 = N687 & N698;
  assign N720 = N687 & yumi_cnt_i[4];
  assign N721 = N689 & N698;
  assign N722 = N689 & yumi_cnt_i[4];
  assign N723 = N691 & N698;
  assign N724 = N691 & yumi_cnt_i[4];
  assign N725 = N693 & N698;
  assign N726 = N693 & yumi_cnt_i[4];
  assign N727 = N695 & N698;
  assign N728 = N695 & yumi_cnt_i[4];
  assign N729 = N697 & N698;
  assign N730 = N697 & yumi_cnt_i[4];
  assign N731 = ~yumi_cnt_i[5];
  assign N732 = N699 & N731;
  assign N733 = N699 & yumi_cnt_i[5];
  assign N734 = N701 & N731;
  assign N735 = N701 & yumi_cnt_i[5];
  assign N736 = N703 & N731;
  assign N737 = N703 & yumi_cnt_i[5];
  assign N738 = N705 & N731;
  assign N739 = N705 & yumi_cnt_i[5];
  assign N740 = N707 & N731;
  assign N741 = N707 & yumi_cnt_i[5];
  assign N742 = N709 & N731;
  assign N743 = N709 & yumi_cnt_i[5];
  assign N744 = N711 & N731;
  assign N745 = N711 & yumi_cnt_i[5];
  assign N746 = N713 & N731;
  assign N747 = N713 & yumi_cnt_i[5];
  assign N748 = N715 & N731;
  assign N749 = N715 & yumi_cnt_i[5];
  assign N750 = N717 & N731;
  assign N751 = N717 & yumi_cnt_i[5];
  assign N752 = N719 & N731;
  assign N753 = N719 & yumi_cnt_i[5];
  assign N754 = N721 & N731;
  assign N755 = N721 & yumi_cnt_i[5];
  assign N756 = N723 & N731;
  assign N757 = N723 & yumi_cnt_i[5];
  assign N758 = N725 & N731;
  assign N759 = N725 & yumi_cnt_i[5];
  assign N760 = N727 & N731;
  assign N761 = N727 & yumi_cnt_i[5];
  assign N762 = N729 & N731;
  assign N763 = N729 & yumi_cnt_i[5];
  assign N764 = N700 & N731;
  assign N765 = N700 & yumi_cnt_i[5];
  assign N766 = N702 & N731;
  assign N767 = N702 & yumi_cnt_i[5];
  assign N768 = N704 & N731;
  assign N769 = N704 & yumi_cnt_i[5];
  assign N770 = N706 & N731;
  assign N771 = N706 & yumi_cnt_i[5];
  assign N772 = N708 & N731;
  assign N773 = N708 & yumi_cnt_i[5];
  assign N774 = N710 & N731;
  assign N775 = N710 & yumi_cnt_i[5];
  assign N776 = N712 & N731;
  assign N777 = N712 & yumi_cnt_i[5];
  assign N778 = N714 & N731;
  assign N779 = N714 & yumi_cnt_i[5];
  assign N780 = N716 & N731;
  assign N781 = N716 & yumi_cnt_i[5];
  assign N782 = N718 & N731;
  assign N783 = N718 & yumi_cnt_i[5];
  assign N784 = N720 & N731;
  assign N785 = N720 & yumi_cnt_i[5];
  assign N786 = N722 & N731;
  assign N787 = N722 & yumi_cnt_i[5];
  assign N788 = N724 & N731;
  assign N789 = N724 & yumi_cnt_i[5];
  assign N790 = N726 & N731;
  assign N791 = N726 & yumi_cnt_i[5];
  assign N792 = N728 & N731;
  assign N793 = N728 & yumi_cnt_i[5];
  assign N794 = N730 & N731;
  assign N795 = N730 & yumi_cnt_i[5];

  always @(posedge clk_i) begin
    if(reset_i) begin
      valid_r_31_sv2v_reg <= 1'b0;
      valid_r_30_sv2v_reg <= 1'b0;
      valid_r_29_sv2v_reg <= 1'b0;
      valid_r_28_sv2v_reg <= 1'b0;
      valid_r_27_sv2v_reg <= 1'b0;
      valid_r_26_sv2v_reg <= 1'b0;
      valid_r_25_sv2v_reg <= 1'b0;
      valid_r_24_sv2v_reg <= 1'b0;
      valid_r_23_sv2v_reg <= 1'b0;
      valid_r_22_sv2v_reg <= 1'b0;
      valid_r_21_sv2v_reg <= 1'b0;
      valid_r_20_sv2v_reg <= 1'b0;
      valid_r_19_sv2v_reg <= 1'b0;
      valid_r_18_sv2v_reg <= 1'b0;
      valid_r_17_sv2v_reg <= 1'b0;
      valid_r_16_sv2v_reg <= 1'b0;
      valid_r_15_sv2v_reg <= 1'b0;
      valid_r_14_sv2v_reg <= 1'b0;
      valid_r_13_sv2v_reg <= 1'b0;
      valid_r_12_sv2v_reg <= 1'b0;
      valid_r_11_sv2v_reg <= 1'b0;
      valid_r_10_sv2v_reg <= 1'b0;
      valid_r_9_sv2v_reg <= 1'b0;
      valid_r_8_sv2v_reg <= 1'b0;
      valid_r_7_sv2v_reg <= 1'b0;
      valid_r_6_sv2v_reg <= 1'b0;
      valid_r_5_sv2v_reg <= 1'b0;
      valid_r_4_sv2v_reg <= 1'b0;
      valid_r_3_sv2v_reg <= 1'b0;
      valid_r_2_sv2v_reg <= 1'b0;
      valid_r_1_sv2v_reg <= 1'b0;
      valid_r_0_sv2v_reg <= 1'b0;
      num_els_r_5_sv2v_reg <= 1'b0;
      num_els_r_4_sv2v_reg <= 1'b0;
      num_els_r_3_sv2v_reg <= 1'b0;
      num_els_r_2_sv2v_reg <= 1'b0;
      num_els_r_1_sv2v_reg <= 1'b0;
      num_els_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      valid_r_31_sv2v_reg <= valid_nn[31];
      valid_r_30_sv2v_reg <= valid_nn[30];
      valid_r_29_sv2v_reg <= valid_nn[29];
      valid_r_28_sv2v_reg <= valid_nn[28];
      valid_r_27_sv2v_reg <= valid_nn[27];
      valid_r_26_sv2v_reg <= valid_nn[26];
      valid_r_25_sv2v_reg <= valid_nn[25];
      valid_r_24_sv2v_reg <= valid_nn[24];
      valid_r_23_sv2v_reg <= valid_nn[23];
      valid_r_22_sv2v_reg <= valid_nn[22];
      valid_r_21_sv2v_reg <= valid_nn[21];
      valid_r_20_sv2v_reg <= valid_nn[20];
      valid_r_19_sv2v_reg <= valid_nn[19];
      valid_r_18_sv2v_reg <= valid_nn[18];
      valid_r_17_sv2v_reg <= valid_nn[17];
      valid_r_16_sv2v_reg <= valid_nn[16];
      valid_r_15_sv2v_reg <= valid_nn[15];
      valid_r_14_sv2v_reg <= valid_nn[14];
      valid_r_13_sv2v_reg <= valid_nn[13];
      valid_r_12_sv2v_reg <= valid_nn[12];
      valid_r_11_sv2v_reg <= valid_nn[11];
      valid_r_10_sv2v_reg <= valid_nn[10];
      valid_r_9_sv2v_reg <= valid_nn[9];
      valid_r_8_sv2v_reg <= valid_nn[8];
      valid_r_7_sv2v_reg <= valid_nn[7];
      valid_r_6_sv2v_reg <= valid_nn[6];
      valid_r_5_sv2v_reg <= valid_nn[5];
      valid_r_4_sv2v_reg <= valid_nn[4];
      valid_r_3_sv2v_reg <= valid_nn[3];
      valid_r_2_sv2v_reg <= valid_nn[2];
      valid_r_1_sv2v_reg <= valid_nn[1];
      valid_r_0_sv2v_reg <= valid_nn[0];
      num_els_r_5_sv2v_reg <= num_els_n[5];
      num_els_r_4_sv2v_reg <= num_els_n[4];
      num_els_r_3_sv2v_reg <= num_els_n[3];
      num_els_r_2_sv2v_reg <= num_els_n[2];
      num_els_r_1_sv2v_reg <= num_els_n[1];
      num_els_r_0_sv2v_reg <= num_els_n[0];
    end 
    if(1'b1) begin
      data_r_511_sv2v_reg <= data_nn[511];
      data_r_510_sv2v_reg <= data_nn[510];
      data_r_509_sv2v_reg <= data_nn[509];
      data_r_508_sv2v_reg <= data_nn[508];
      data_r_507_sv2v_reg <= data_nn[507];
      data_r_506_sv2v_reg <= data_nn[506];
      data_r_505_sv2v_reg <= data_nn[505];
      data_r_504_sv2v_reg <= data_nn[504];
      data_r_503_sv2v_reg <= data_nn[503];
      data_r_502_sv2v_reg <= data_nn[502];
      data_r_501_sv2v_reg <= data_nn[501];
      data_r_500_sv2v_reg <= data_nn[500];
      data_r_499_sv2v_reg <= data_nn[499];
      data_r_498_sv2v_reg <= data_nn[498];
      data_r_497_sv2v_reg <= data_nn[497];
      data_r_496_sv2v_reg <= data_nn[496];
      data_r_495_sv2v_reg <= data_nn[495];
      data_r_494_sv2v_reg <= data_nn[494];
      data_r_493_sv2v_reg <= data_nn[493];
      data_r_492_sv2v_reg <= data_nn[492];
      data_r_491_sv2v_reg <= data_nn[491];
      data_r_490_sv2v_reg <= data_nn[490];
      data_r_489_sv2v_reg <= data_nn[489];
      data_r_488_sv2v_reg <= data_nn[488];
      data_r_487_sv2v_reg <= data_nn[487];
      data_r_486_sv2v_reg <= data_nn[486];
      data_r_485_sv2v_reg <= data_nn[485];
      data_r_484_sv2v_reg <= data_nn[484];
      data_r_483_sv2v_reg <= data_nn[483];
      data_r_482_sv2v_reg <= data_nn[482];
      data_r_481_sv2v_reg <= data_nn[481];
      data_r_480_sv2v_reg <= data_nn[480];
      data_r_479_sv2v_reg <= data_nn[479];
      data_r_478_sv2v_reg <= data_nn[478];
      data_r_477_sv2v_reg <= data_nn[477];
      data_r_476_sv2v_reg <= data_nn[476];
      data_r_475_sv2v_reg <= data_nn[475];
      data_r_474_sv2v_reg <= data_nn[474];
      data_r_473_sv2v_reg <= data_nn[473];
      data_r_472_sv2v_reg <= data_nn[472];
      data_r_471_sv2v_reg <= data_nn[471];
      data_r_470_sv2v_reg <= data_nn[470];
      data_r_469_sv2v_reg <= data_nn[469];
      data_r_468_sv2v_reg <= data_nn[468];
      data_r_467_sv2v_reg <= data_nn[467];
      data_r_466_sv2v_reg <= data_nn[466];
      data_r_465_sv2v_reg <= data_nn[465];
      data_r_464_sv2v_reg <= data_nn[464];
      data_r_463_sv2v_reg <= data_nn[463];
      data_r_462_sv2v_reg <= data_nn[462];
      data_r_461_sv2v_reg <= data_nn[461];
      data_r_460_sv2v_reg <= data_nn[460];
      data_r_459_sv2v_reg <= data_nn[459];
      data_r_458_sv2v_reg <= data_nn[458];
      data_r_457_sv2v_reg <= data_nn[457];
      data_r_456_sv2v_reg <= data_nn[456];
      data_r_455_sv2v_reg <= data_nn[455];
      data_r_454_sv2v_reg <= data_nn[454];
      data_r_453_sv2v_reg <= data_nn[453];
      data_r_452_sv2v_reg <= data_nn[452];
      data_r_451_sv2v_reg <= data_nn[451];
      data_r_450_sv2v_reg <= data_nn[450];
      data_r_449_sv2v_reg <= data_nn[449];
      data_r_448_sv2v_reg <= data_nn[448];
      data_r_447_sv2v_reg <= data_nn[447];
      data_r_446_sv2v_reg <= data_nn[446];
      data_r_445_sv2v_reg <= data_nn[445];
      data_r_444_sv2v_reg <= data_nn[444];
      data_r_443_sv2v_reg <= data_nn[443];
      data_r_442_sv2v_reg <= data_nn[442];
      data_r_441_sv2v_reg <= data_nn[441];
      data_r_440_sv2v_reg <= data_nn[440];
      data_r_439_sv2v_reg <= data_nn[439];
      data_r_438_sv2v_reg <= data_nn[438];
      data_r_437_sv2v_reg <= data_nn[437];
      data_r_436_sv2v_reg <= data_nn[436];
      data_r_435_sv2v_reg <= data_nn[435];
      data_r_434_sv2v_reg <= data_nn[434];
      data_r_433_sv2v_reg <= data_nn[433];
      data_r_432_sv2v_reg <= data_nn[432];
      data_r_431_sv2v_reg <= data_nn[431];
      data_r_430_sv2v_reg <= data_nn[430];
      data_r_429_sv2v_reg <= data_nn[429];
      data_r_428_sv2v_reg <= data_nn[428];
      data_r_427_sv2v_reg <= data_nn[427];
      data_r_426_sv2v_reg <= data_nn[426];
      data_r_425_sv2v_reg <= data_nn[425];
      data_r_424_sv2v_reg <= data_nn[424];
      data_r_423_sv2v_reg <= data_nn[423];
      data_r_422_sv2v_reg <= data_nn[422];
      data_r_421_sv2v_reg <= data_nn[421];
      data_r_420_sv2v_reg <= data_nn[420];
      data_r_419_sv2v_reg <= data_nn[419];
      data_r_418_sv2v_reg <= data_nn[418];
      data_r_417_sv2v_reg <= data_nn[417];
      data_r_416_sv2v_reg <= data_nn[416];
      data_r_415_sv2v_reg <= data_nn[415];
      data_r_414_sv2v_reg <= data_nn[414];
      data_r_413_sv2v_reg <= data_nn[413];
      data_r_412_sv2v_reg <= data_nn[412];
      data_r_411_sv2v_reg <= data_nn[411];
      data_r_410_sv2v_reg <= data_nn[410];
      data_r_409_sv2v_reg <= data_nn[409];
      data_r_408_sv2v_reg <= data_nn[408];
      data_r_407_sv2v_reg <= data_nn[407];
      data_r_406_sv2v_reg <= data_nn[406];
      data_r_405_sv2v_reg <= data_nn[405];
      data_r_404_sv2v_reg <= data_nn[404];
      data_r_403_sv2v_reg <= data_nn[403];
      data_r_402_sv2v_reg <= data_nn[402];
      data_r_401_sv2v_reg <= data_nn[401];
      data_r_400_sv2v_reg <= data_nn[400];
      data_r_399_sv2v_reg <= data_nn[399];
      data_r_398_sv2v_reg <= data_nn[398];
      data_r_397_sv2v_reg <= data_nn[397];
      data_r_396_sv2v_reg <= data_nn[396];
      data_r_395_sv2v_reg <= data_nn[395];
      data_r_394_sv2v_reg <= data_nn[394];
      data_r_393_sv2v_reg <= data_nn[393];
      data_r_392_sv2v_reg <= data_nn[392];
      data_r_391_sv2v_reg <= data_nn[391];
      data_r_390_sv2v_reg <= data_nn[390];
      data_r_389_sv2v_reg <= data_nn[389];
      data_r_388_sv2v_reg <= data_nn[388];
      data_r_387_sv2v_reg <= data_nn[387];
      data_r_386_sv2v_reg <= data_nn[386];
      data_r_385_sv2v_reg <= data_nn[385];
      data_r_384_sv2v_reg <= data_nn[384];
      data_r_383_sv2v_reg <= data_nn[383];
      data_r_382_sv2v_reg <= data_nn[382];
      data_r_381_sv2v_reg <= data_nn[381];
      data_r_380_sv2v_reg <= data_nn[380];
      data_r_379_sv2v_reg <= data_nn[379];
      data_r_378_sv2v_reg <= data_nn[378];
      data_r_377_sv2v_reg <= data_nn[377];
      data_r_376_sv2v_reg <= data_nn[376];
      data_r_375_sv2v_reg <= data_nn[375];
      data_r_374_sv2v_reg <= data_nn[374];
      data_r_373_sv2v_reg <= data_nn[373];
      data_r_372_sv2v_reg <= data_nn[372];
      data_r_371_sv2v_reg <= data_nn[371];
      data_r_370_sv2v_reg <= data_nn[370];
      data_r_369_sv2v_reg <= data_nn[369];
      data_r_368_sv2v_reg <= data_nn[368];
      data_r_367_sv2v_reg <= data_nn[367];
      data_r_366_sv2v_reg <= data_nn[366];
      data_r_365_sv2v_reg <= data_nn[365];
      data_r_364_sv2v_reg <= data_nn[364];
      data_r_363_sv2v_reg <= data_nn[363];
      data_r_362_sv2v_reg <= data_nn[362];
      data_r_361_sv2v_reg <= data_nn[361];
      data_r_360_sv2v_reg <= data_nn[360];
      data_r_359_sv2v_reg <= data_nn[359];
      data_r_358_sv2v_reg <= data_nn[358];
      data_r_357_sv2v_reg <= data_nn[357];
      data_r_356_sv2v_reg <= data_nn[356];
      data_r_355_sv2v_reg <= data_nn[355];
      data_r_354_sv2v_reg <= data_nn[354];
      data_r_353_sv2v_reg <= data_nn[353];
      data_r_352_sv2v_reg <= data_nn[352];
      data_r_351_sv2v_reg <= data_nn[351];
      data_r_350_sv2v_reg <= data_nn[350];
      data_r_349_sv2v_reg <= data_nn[349];
      data_r_348_sv2v_reg <= data_nn[348];
      data_r_347_sv2v_reg <= data_nn[347];
      data_r_346_sv2v_reg <= data_nn[346];
      data_r_345_sv2v_reg <= data_nn[345];
      data_r_344_sv2v_reg <= data_nn[344];
      data_r_343_sv2v_reg <= data_nn[343];
      data_r_342_sv2v_reg <= data_nn[342];
      data_r_341_sv2v_reg <= data_nn[341];
      data_r_340_sv2v_reg <= data_nn[340];
      data_r_339_sv2v_reg <= data_nn[339];
      data_r_338_sv2v_reg <= data_nn[338];
      data_r_337_sv2v_reg <= data_nn[337];
      data_r_336_sv2v_reg <= data_nn[336];
      data_r_335_sv2v_reg <= data_nn[335];
      data_r_334_sv2v_reg <= data_nn[334];
      data_r_333_sv2v_reg <= data_nn[333];
      data_r_332_sv2v_reg <= data_nn[332];
      data_r_331_sv2v_reg <= data_nn[331];
      data_r_330_sv2v_reg <= data_nn[330];
      data_r_329_sv2v_reg <= data_nn[329];
      data_r_328_sv2v_reg <= data_nn[328];
      data_r_327_sv2v_reg <= data_nn[327];
      data_r_326_sv2v_reg <= data_nn[326];
      data_r_325_sv2v_reg <= data_nn[325];
      data_r_324_sv2v_reg <= data_nn[324];
      data_r_323_sv2v_reg <= data_nn[323];
      data_r_322_sv2v_reg <= data_nn[322];
      data_r_321_sv2v_reg <= data_nn[321];
      data_r_320_sv2v_reg <= data_nn[320];
      data_r_319_sv2v_reg <= data_nn[319];
      data_r_318_sv2v_reg <= data_nn[318];
      data_r_317_sv2v_reg <= data_nn[317];
      data_r_316_sv2v_reg <= data_nn[316];
      data_r_315_sv2v_reg <= data_nn[315];
      data_r_314_sv2v_reg <= data_nn[314];
      data_r_313_sv2v_reg <= data_nn[313];
      data_r_312_sv2v_reg <= data_nn[312];
      data_r_311_sv2v_reg <= data_nn[311];
      data_r_310_sv2v_reg <= data_nn[310];
      data_r_309_sv2v_reg <= data_nn[309];
      data_r_308_sv2v_reg <= data_nn[308];
      data_r_307_sv2v_reg <= data_nn[307];
      data_r_306_sv2v_reg <= data_nn[306];
      data_r_305_sv2v_reg <= data_nn[305];
      data_r_304_sv2v_reg <= data_nn[304];
      data_r_303_sv2v_reg <= data_nn[303];
      data_r_302_sv2v_reg <= data_nn[302];
      data_r_301_sv2v_reg <= data_nn[301];
      data_r_300_sv2v_reg <= data_nn[300];
      data_r_299_sv2v_reg <= data_nn[299];
      data_r_298_sv2v_reg <= data_nn[298];
      data_r_297_sv2v_reg <= data_nn[297];
      data_r_296_sv2v_reg <= data_nn[296];
      data_r_295_sv2v_reg <= data_nn[295];
      data_r_294_sv2v_reg <= data_nn[294];
      data_r_293_sv2v_reg <= data_nn[293];
      data_r_292_sv2v_reg <= data_nn[292];
      data_r_291_sv2v_reg <= data_nn[291];
      data_r_290_sv2v_reg <= data_nn[290];
      data_r_289_sv2v_reg <= data_nn[289];
      data_r_288_sv2v_reg <= data_nn[288];
      data_r_287_sv2v_reg <= data_nn[287];
      data_r_286_sv2v_reg <= data_nn[286];
      data_r_285_sv2v_reg <= data_nn[285];
      data_r_284_sv2v_reg <= data_nn[284];
      data_r_283_sv2v_reg <= data_nn[283];
      data_r_282_sv2v_reg <= data_nn[282];
      data_r_281_sv2v_reg <= data_nn[281];
      data_r_280_sv2v_reg <= data_nn[280];
      data_r_279_sv2v_reg <= data_nn[279];
      data_r_278_sv2v_reg <= data_nn[278];
      data_r_277_sv2v_reg <= data_nn[277];
      data_r_276_sv2v_reg <= data_nn[276];
      data_r_275_sv2v_reg <= data_nn[275];
      data_r_274_sv2v_reg <= data_nn[274];
      data_r_273_sv2v_reg <= data_nn[273];
      data_r_272_sv2v_reg <= data_nn[272];
      data_r_271_sv2v_reg <= data_nn[271];
      data_r_270_sv2v_reg <= data_nn[270];
      data_r_269_sv2v_reg <= data_nn[269];
      data_r_268_sv2v_reg <= data_nn[268];
      data_r_267_sv2v_reg <= data_nn[267];
      data_r_266_sv2v_reg <= data_nn[266];
      data_r_265_sv2v_reg <= data_nn[265];
      data_r_264_sv2v_reg <= data_nn[264];
      data_r_263_sv2v_reg <= data_nn[263];
      data_r_262_sv2v_reg <= data_nn[262];
      data_r_261_sv2v_reg <= data_nn[261];
      data_r_260_sv2v_reg <= data_nn[260];
      data_r_259_sv2v_reg <= data_nn[259];
      data_r_258_sv2v_reg <= data_nn[258];
      data_r_257_sv2v_reg <= data_nn[257];
      data_r_256_sv2v_reg <= data_nn[256];
      data_r_255_sv2v_reg <= data_nn[255];
      data_r_254_sv2v_reg <= data_nn[254];
      data_r_253_sv2v_reg <= data_nn[253];
      data_r_252_sv2v_reg <= data_nn[252];
      data_r_251_sv2v_reg <= data_nn[251];
      data_r_250_sv2v_reg <= data_nn[250];
      data_r_249_sv2v_reg <= data_nn[249];
      data_r_248_sv2v_reg <= data_nn[248];
      data_r_247_sv2v_reg <= data_nn[247];
      data_r_246_sv2v_reg <= data_nn[246];
      data_r_245_sv2v_reg <= data_nn[245];
      data_r_244_sv2v_reg <= data_nn[244];
      data_r_243_sv2v_reg <= data_nn[243];
      data_r_242_sv2v_reg <= data_nn[242];
      data_r_241_sv2v_reg <= data_nn[241];
      data_r_240_sv2v_reg <= data_nn[240];
      data_r_239_sv2v_reg <= data_nn[239];
      data_r_238_sv2v_reg <= data_nn[238];
      data_r_237_sv2v_reg <= data_nn[237];
      data_r_236_sv2v_reg <= data_nn[236];
      data_r_235_sv2v_reg <= data_nn[235];
      data_r_234_sv2v_reg <= data_nn[234];
      data_r_233_sv2v_reg <= data_nn[233];
      data_r_232_sv2v_reg <= data_nn[232];
      data_r_231_sv2v_reg <= data_nn[231];
      data_r_230_sv2v_reg <= data_nn[230];
      data_r_229_sv2v_reg <= data_nn[229];
      data_r_228_sv2v_reg <= data_nn[228];
      data_r_227_sv2v_reg <= data_nn[227];
      data_r_226_sv2v_reg <= data_nn[226];
      data_r_225_sv2v_reg <= data_nn[225];
      data_r_224_sv2v_reg <= data_nn[224];
      data_r_223_sv2v_reg <= data_nn[223];
      data_r_222_sv2v_reg <= data_nn[222];
      data_r_221_sv2v_reg <= data_nn[221];
      data_r_220_sv2v_reg <= data_nn[220];
      data_r_219_sv2v_reg <= data_nn[219];
      data_r_218_sv2v_reg <= data_nn[218];
      data_r_217_sv2v_reg <= data_nn[217];
      data_r_216_sv2v_reg <= data_nn[216];
      data_r_215_sv2v_reg <= data_nn[215];
      data_r_214_sv2v_reg <= data_nn[214];
      data_r_213_sv2v_reg <= data_nn[213];
      data_r_212_sv2v_reg <= data_nn[212];
      data_r_211_sv2v_reg <= data_nn[211];
      data_r_210_sv2v_reg <= data_nn[210];
      data_r_209_sv2v_reg <= data_nn[209];
      data_r_208_sv2v_reg <= data_nn[208];
      data_r_207_sv2v_reg <= data_nn[207];
      data_r_206_sv2v_reg <= data_nn[206];
      data_r_205_sv2v_reg <= data_nn[205];
      data_r_204_sv2v_reg <= data_nn[204];
      data_r_203_sv2v_reg <= data_nn[203];
      data_r_202_sv2v_reg <= data_nn[202];
      data_r_201_sv2v_reg <= data_nn[201];
      data_r_200_sv2v_reg <= data_nn[200];
      data_r_199_sv2v_reg <= data_nn[199];
      data_r_198_sv2v_reg <= data_nn[198];
      data_r_197_sv2v_reg <= data_nn[197];
      data_r_196_sv2v_reg <= data_nn[196];
      data_r_195_sv2v_reg <= data_nn[195];
      data_r_194_sv2v_reg <= data_nn[194];
      data_r_193_sv2v_reg <= data_nn[193];
      data_r_192_sv2v_reg <= data_nn[192];
      data_r_191_sv2v_reg <= data_nn[191];
      data_r_190_sv2v_reg <= data_nn[190];
      data_r_189_sv2v_reg <= data_nn[189];
      data_r_188_sv2v_reg <= data_nn[188];
      data_r_187_sv2v_reg <= data_nn[187];
      data_r_186_sv2v_reg <= data_nn[186];
      data_r_185_sv2v_reg <= data_nn[185];
      data_r_184_sv2v_reg <= data_nn[184];
      data_r_183_sv2v_reg <= data_nn[183];
      data_r_182_sv2v_reg <= data_nn[182];
      data_r_181_sv2v_reg <= data_nn[181];
      data_r_180_sv2v_reg <= data_nn[180];
      data_r_179_sv2v_reg <= data_nn[179];
      data_r_178_sv2v_reg <= data_nn[178];
      data_r_177_sv2v_reg <= data_nn[177];
      data_r_176_sv2v_reg <= data_nn[176];
      data_r_175_sv2v_reg <= data_nn[175];
      data_r_174_sv2v_reg <= data_nn[174];
      data_r_173_sv2v_reg <= data_nn[173];
      data_r_172_sv2v_reg <= data_nn[172];
      data_r_171_sv2v_reg <= data_nn[171];
      data_r_170_sv2v_reg <= data_nn[170];
      data_r_169_sv2v_reg <= data_nn[169];
      data_r_168_sv2v_reg <= data_nn[168];
      data_r_167_sv2v_reg <= data_nn[167];
      data_r_166_sv2v_reg <= data_nn[166];
      data_r_165_sv2v_reg <= data_nn[165];
      data_r_164_sv2v_reg <= data_nn[164];
      data_r_163_sv2v_reg <= data_nn[163];
      data_r_162_sv2v_reg <= data_nn[162];
      data_r_161_sv2v_reg <= data_nn[161];
      data_r_160_sv2v_reg <= data_nn[160];
      data_r_159_sv2v_reg <= data_nn[159];
      data_r_158_sv2v_reg <= data_nn[158];
      data_r_157_sv2v_reg <= data_nn[157];
      data_r_156_sv2v_reg <= data_nn[156];
      data_r_155_sv2v_reg <= data_nn[155];
      data_r_154_sv2v_reg <= data_nn[154];
      data_r_153_sv2v_reg <= data_nn[153];
      data_r_152_sv2v_reg <= data_nn[152];
      data_r_151_sv2v_reg <= data_nn[151];
      data_r_150_sv2v_reg <= data_nn[150];
      data_r_149_sv2v_reg <= data_nn[149];
      data_r_148_sv2v_reg <= data_nn[148];
      data_r_147_sv2v_reg <= data_nn[147];
      data_r_146_sv2v_reg <= data_nn[146];
      data_r_145_sv2v_reg <= data_nn[145];
      data_r_144_sv2v_reg <= data_nn[144];
      data_r_143_sv2v_reg <= data_nn[143];
      data_r_142_sv2v_reg <= data_nn[142];
      data_r_141_sv2v_reg <= data_nn[141];
      data_r_140_sv2v_reg <= data_nn[140];
      data_r_139_sv2v_reg <= data_nn[139];
      data_r_138_sv2v_reg <= data_nn[138];
      data_r_137_sv2v_reg <= data_nn[137];
      data_r_136_sv2v_reg <= data_nn[136];
      data_r_135_sv2v_reg <= data_nn[135];
      data_r_134_sv2v_reg <= data_nn[134];
      data_r_133_sv2v_reg <= data_nn[133];
      data_r_132_sv2v_reg <= data_nn[132];
      data_r_131_sv2v_reg <= data_nn[131];
      data_r_130_sv2v_reg <= data_nn[130];
      data_r_129_sv2v_reg <= data_nn[129];
      data_r_128_sv2v_reg <= data_nn[128];
      data_r_127_sv2v_reg <= data_nn[127];
      data_r_126_sv2v_reg <= data_nn[126];
      data_r_125_sv2v_reg <= data_nn[125];
      data_r_124_sv2v_reg <= data_nn[124];
      data_r_123_sv2v_reg <= data_nn[123];
      data_r_122_sv2v_reg <= data_nn[122];
      data_r_121_sv2v_reg <= data_nn[121];
      data_r_120_sv2v_reg <= data_nn[120];
      data_r_119_sv2v_reg <= data_nn[119];
      data_r_118_sv2v_reg <= data_nn[118];
      data_r_117_sv2v_reg <= data_nn[117];
      data_r_116_sv2v_reg <= data_nn[116];
      data_r_115_sv2v_reg <= data_nn[115];
      data_r_114_sv2v_reg <= data_nn[114];
      data_r_113_sv2v_reg <= data_nn[113];
      data_r_112_sv2v_reg <= data_nn[112];
      data_r_111_sv2v_reg <= data_nn[111];
      data_r_110_sv2v_reg <= data_nn[110];
      data_r_109_sv2v_reg <= data_nn[109];
      data_r_108_sv2v_reg <= data_nn[108];
      data_r_107_sv2v_reg <= data_nn[107];
      data_r_106_sv2v_reg <= data_nn[106];
      data_r_105_sv2v_reg <= data_nn[105];
      data_r_104_sv2v_reg <= data_nn[104];
      data_r_103_sv2v_reg <= data_nn[103];
      data_r_102_sv2v_reg <= data_nn[102];
      data_r_101_sv2v_reg <= data_nn[101];
      data_r_100_sv2v_reg <= data_nn[100];
      data_r_99_sv2v_reg <= data_nn[99];
      data_r_98_sv2v_reg <= data_nn[98];
      data_r_97_sv2v_reg <= data_nn[97];
      data_r_96_sv2v_reg <= data_nn[96];
      data_r_95_sv2v_reg <= data_nn[95];
      data_r_94_sv2v_reg <= data_nn[94];
      data_r_93_sv2v_reg <= data_nn[93];
      data_r_92_sv2v_reg <= data_nn[92];
      data_r_91_sv2v_reg <= data_nn[91];
      data_r_90_sv2v_reg <= data_nn[90];
      data_r_89_sv2v_reg <= data_nn[89];
      data_r_88_sv2v_reg <= data_nn[88];
      data_r_87_sv2v_reg <= data_nn[87];
      data_r_86_sv2v_reg <= data_nn[86];
      data_r_85_sv2v_reg <= data_nn[85];
      data_r_84_sv2v_reg <= data_nn[84];
      data_r_83_sv2v_reg <= data_nn[83];
      data_r_82_sv2v_reg <= data_nn[82];
      data_r_81_sv2v_reg <= data_nn[81];
      data_r_80_sv2v_reg <= data_nn[80];
      data_r_79_sv2v_reg <= data_nn[79];
      data_r_78_sv2v_reg <= data_nn[78];
      data_r_77_sv2v_reg <= data_nn[77];
      data_r_76_sv2v_reg <= data_nn[76];
      data_r_75_sv2v_reg <= data_nn[75];
      data_r_74_sv2v_reg <= data_nn[74];
      data_r_73_sv2v_reg <= data_nn[73];
      data_r_72_sv2v_reg <= data_nn[72];
      data_r_71_sv2v_reg <= data_nn[71];
      data_r_70_sv2v_reg <= data_nn[70];
      data_r_69_sv2v_reg <= data_nn[69];
      data_r_68_sv2v_reg <= data_nn[68];
      data_r_67_sv2v_reg <= data_nn[67];
      data_r_66_sv2v_reg <= data_nn[66];
      data_r_65_sv2v_reg <= data_nn[65];
      data_r_64_sv2v_reg <= data_nn[64];
      data_r_63_sv2v_reg <= data_nn[63];
      data_r_62_sv2v_reg <= data_nn[62];
      data_r_61_sv2v_reg <= data_nn[61];
      data_r_60_sv2v_reg <= data_nn[60];
      data_r_59_sv2v_reg <= data_nn[59];
      data_r_58_sv2v_reg <= data_nn[58];
      data_r_57_sv2v_reg <= data_nn[57];
      data_r_56_sv2v_reg <= data_nn[56];
      data_r_55_sv2v_reg <= data_nn[55];
      data_r_54_sv2v_reg <= data_nn[54];
      data_r_53_sv2v_reg <= data_nn[53];
      data_r_52_sv2v_reg <= data_nn[52];
      data_r_51_sv2v_reg <= data_nn[51];
      data_r_50_sv2v_reg <= data_nn[50];
      data_r_49_sv2v_reg <= data_nn[49];
      data_r_48_sv2v_reg <= data_nn[48];
      data_r_47_sv2v_reg <= data_nn[47];
      data_r_46_sv2v_reg <= data_nn[46];
      data_r_45_sv2v_reg <= data_nn[45];
      data_r_44_sv2v_reg <= data_nn[44];
      data_r_43_sv2v_reg <= data_nn[43];
      data_r_42_sv2v_reg <= data_nn[42];
      data_r_41_sv2v_reg <= data_nn[41];
      data_r_40_sv2v_reg <= data_nn[40];
      data_r_39_sv2v_reg <= data_nn[39];
      data_r_38_sv2v_reg <= data_nn[38];
      data_r_37_sv2v_reg <= data_nn[37];
      data_r_36_sv2v_reg <= data_nn[36];
      data_r_35_sv2v_reg <= data_nn[35];
      data_r_34_sv2v_reg <= data_nn[34];
      data_r_33_sv2v_reg <= data_nn[33];
      data_r_32_sv2v_reg <= data_nn[32];
      data_r_31_sv2v_reg <= data_nn[31];
      data_r_30_sv2v_reg <= data_nn[30];
      data_r_29_sv2v_reg <= data_nn[29];
      data_r_28_sv2v_reg <= data_nn[28];
      data_r_27_sv2v_reg <= data_nn[27];
      data_r_26_sv2v_reg <= data_nn[26];
      data_r_25_sv2v_reg <= data_nn[25];
      data_r_24_sv2v_reg <= data_nn[24];
      data_r_23_sv2v_reg <= data_nn[23];
      data_r_22_sv2v_reg <= data_nn[22];
      data_r_21_sv2v_reg <= data_nn[21];
      data_r_20_sv2v_reg <= data_nn[20];
      data_r_19_sv2v_reg <= data_nn[19];
      data_r_18_sv2v_reg <= data_nn[18];
      data_r_17_sv2v_reg <= data_nn[17];
      data_r_16_sv2v_reg <= data_nn[16];
      data_r_15_sv2v_reg <= data_nn[15];
      data_r_14_sv2v_reg <= data_nn[14];
      data_r_13_sv2v_reg <= data_nn[13];
      data_r_12_sv2v_reg <= data_nn[12];
      data_r_11_sv2v_reg <= data_nn[11];
      data_r_10_sv2v_reg <= data_nn[10];
      data_r_9_sv2v_reg <= data_nn[9];
      data_r_8_sv2v_reg <= data_nn[8];
      data_r_7_sv2v_reg <= data_nn[7];
      data_r_6_sv2v_reg <= data_nn[6];
      data_r_5_sv2v_reg <= data_nn[5];
      data_r_4_sv2v_reg <= data_nn[4];
      data_r_3_sv2v_reg <= data_nn[3];
      data_r_2_sv2v_reg <= data_nn[2];
      data_r_1_sv2v_reg <= data_nn[1];
      data_r_0_sv2v_reg <= data_nn[0];
    end 
  end


endmodule

