module top(output int o);
   shortreal a = 0.5;
   assign o = int'(2 * a);
endmodule
