module top(output logic[7:0] o);
   assign o = '{default: 1};
endmodule
