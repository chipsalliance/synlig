module top(output int o);
   parameter int P = 1;
   assign o = P + 2;
endmodule
