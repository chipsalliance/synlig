package my_pkg;
   parameter int A__B = 1;
endpackage // my_pkg
