

module top
(
  i,
  o
);

  input [255:0] i;
  output [255:0] o;

  bsg_transpose
  wrapper
  (
    .i(i),
    .o(o)
  );


endmodule



module bsg_transpose
(
  i,
  o
);

  input [255:0] i;
  output [255:0] o;
  wire [255:0] o;
  assign o[255] = i[255];
  assign o[254] = i[239];
  assign o[253] = i[223];
  assign o[252] = i[207];
  assign o[251] = i[191];
  assign o[250] = i[175];
  assign o[249] = i[159];
  assign o[248] = i[143];
  assign o[247] = i[127];
  assign o[246] = i[111];
  assign o[245] = i[95];
  assign o[244] = i[79];
  assign o[243] = i[63];
  assign o[242] = i[47];
  assign o[241] = i[31];
  assign o[240] = i[15];
  assign o[239] = i[254];
  assign o[238] = i[238];
  assign o[237] = i[222];
  assign o[236] = i[206];
  assign o[235] = i[190];
  assign o[234] = i[174];
  assign o[233] = i[158];
  assign o[232] = i[142];
  assign o[231] = i[126];
  assign o[230] = i[110];
  assign o[229] = i[94];
  assign o[228] = i[78];
  assign o[227] = i[62];
  assign o[226] = i[46];
  assign o[225] = i[30];
  assign o[224] = i[14];
  assign o[223] = i[253];
  assign o[222] = i[237];
  assign o[221] = i[221];
  assign o[220] = i[205];
  assign o[219] = i[189];
  assign o[218] = i[173];
  assign o[217] = i[157];
  assign o[216] = i[141];
  assign o[215] = i[125];
  assign o[214] = i[109];
  assign o[213] = i[93];
  assign o[212] = i[77];
  assign o[211] = i[61];
  assign o[210] = i[45];
  assign o[209] = i[29];
  assign o[208] = i[13];
  assign o[207] = i[252];
  assign o[206] = i[236];
  assign o[205] = i[220];
  assign o[204] = i[204];
  assign o[203] = i[188];
  assign o[202] = i[172];
  assign o[201] = i[156];
  assign o[200] = i[140];
  assign o[199] = i[124];
  assign o[198] = i[108];
  assign o[197] = i[92];
  assign o[196] = i[76];
  assign o[195] = i[60];
  assign o[194] = i[44];
  assign o[193] = i[28];
  assign o[192] = i[12];
  assign o[191] = i[251];
  assign o[190] = i[235];
  assign o[189] = i[219];
  assign o[188] = i[203];
  assign o[187] = i[187];
  assign o[186] = i[171];
  assign o[185] = i[155];
  assign o[184] = i[139];
  assign o[183] = i[123];
  assign o[182] = i[107];
  assign o[181] = i[91];
  assign o[180] = i[75];
  assign o[179] = i[59];
  assign o[178] = i[43];
  assign o[177] = i[27];
  assign o[176] = i[11];
  assign o[175] = i[250];
  assign o[174] = i[234];
  assign o[173] = i[218];
  assign o[172] = i[202];
  assign o[171] = i[186];
  assign o[170] = i[170];
  assign o[169] = i[154];
  assign o[168] = i[138];
  assign o[167] = i[122];
  assign o[166] = i[106];
  assign o[165] = i[90];
  assign o[164] = i[74];
  assign o[163] = i[58];
  assign o[162] = i[42];
  assign o[161] = i[26];
  assign o[160] = i[10];
  assign o[159] = i[249];
  assign o[158] = i[233];
  assign o[157] = i[217];
  assign o[156] = i[201];
  assign o[155] = i[185];
  assign o[154] = i[169];
  assign o[153] = i[153];
  assign o[152] = i[137];
  assign o[151] = i[121];
  assign o[150] = i[105];
  assign o[149] = i[89];
  assign o[148] = i[73];
  assign o[147] = i[57];
  assign o[146] = i[41];
  assign o[145] = i[25];
  assign o[144] = i[9];
  assign o[143] = i[248];
  assign o[142] = i[232];
  assign o[141] = i[216];
  assign o[140] = i[200];
  assign o[139] = i[184];
  assign o[138] = i[168];
  assign o[137] = i[152];
  assign o[136] = i[136];
  assign o[135] = i[120];
  assign o[134] = i[104];
  assign o[133] = i[88];
  assign o[132] = i[72];
  assign o[131] = i[56];
  assign o[130] = i[40];
  assign o[129] = i[24];
  assign o[128] = i[8];
  assign o[127] = i[247];
  assign o[126] = i[231];
  assign o[125] = i[215];
  assign o[124] = i[199];
  assign o[123] = i[183];
  assign o[122] = i[167];
  assign o[121] = i[151];
  assign o[120] = i[135];
  assign o[119] = i[119];
  assign o[118] = i[103];
  assign o[117] = i[87];
  assign o[116] = i[71];
  assign o[115] = i[55];
  assign o[114] = i[39];
  assign o[113] = i[23];
  assign o[112] = i[7];
  assign o[111] = i[246];
  assign o[110] = i[230];
  assign o[109] = i[214];
  assign o[108] = i[198];
  assign o[107] = i[182];
  assign o[106] = i[166];
  assign o[105] = i[150];
  assign o[104] = i[134];
  assign o[103] = i[118];
  assign o[102] = i[102];
  assign o[101] = i[86];
  assign o[100] = i[70];
  assign o[99] = i[54];
  assign o[98] = i[38];
  assign o[97] = i[22];
  assign o[96] = i[6];
  assign o[95] = i[245];
  assign o[94] = i[229];
  assign o[93] = i[213];
  assign o[92] = i[197];
  assign o[91] = i[181];
  assign o[90] = i[165];
  assign o[89] = i[149];
  assign o[88] = i[133];
  assign o[87] = i[117];
  assign o[86] = i[101];
  assign o[85] = i[85];
  assign o[84] = i[69];
  assign o[83] = i[53];
  assign o[82] = i[37];
  assign o[81] = i[21];
  assign o[80] = i[5];
  assign o[79] = i[244];
  assign o[78] = i[228];
  assign o[77] = i[212];
  assign o[76] = i[196];
  assign o[75] = i[180];
  assign o[74] = i[164];
  assign o[73] = i[148];
  assign o[72] = i[132];
  assign o[71] = i[116];
  assign o[70] = i[100];
  assign o[69] = i[84];
  assign o[68] = i[68];
  assign o[67] = i[52];
  assign o[66] = i[36];
  assign o[65] = i[20];
  assign o[64] = i[4];
  assign o[63] = i[243];
  assign o[62] = i[227];
  assign o[61] = i[211];
  assign o[60] = i[195];
  assign o[59] = i[179];
  assign o[58] = i[163];
  assign o[57] = i[147];
  assign o[56] = i[131];
  assign o[55] = i[115];
  assign o[54] = i[99];
  assign o[53] = i[83];
  assign o[52] = i[67];
  assign o[51] = i[51];
  assign o[50] = i[35];
  assign o[49] = i[19];
  assign o[48] = i[3];
  assign o[47] = i[242];
  assign o[46] = i[226];
  assign o[45] = i[210];
  assign o[44] = i[194];
  assign o[43] = i[178];
  assign o[42] = i[162];
  assign o[41] = i[146];
  assign o[40] = i[130];
  assign o[39] = i[114];
  assign o[38] = i[98];
  assign o[37] = i[82];
  assign o[36] = i[66];
  assign o[35] = i[50];
  assign o[34] = i[34];
  assign o[33] = i[18];
  assign o[32] = i[2];
  assign o[31] = i[241];
  assign o[30] = i[225];
  assign o[29] = i[209];
  assign o[28] = i[193];
  assign o[27] = i[177];
  assign o[26] = i[161];
  assign o[25] = i[145];
  assign o[24] = i[129];
  assign o[23] = i[113];
  assign o[22] = i[97];
  assign o[21] = i[81];
  assign o[20] = i[65];
  assign o[19] = i[49];
  assign o[18] = i[33];
  assign o[17] = i[17];
  assign o[16] = i[1];
  assign o[15] = i[240];
  assign o[14] = i[224];
  assign o[13] = i[208];
  assign o[12] = i[192];
  assign o[11] = i[176];
  assign o[10] = i[160];
  assign o[9] = i[144];
  assign o[8] = i[128];
  assign o[7] = i[112];
  assign o[6] = i[96];
  assign o[5] = i[80];
  assign o[4] = i[64];
  assign o[3] = i[48];
  assign o[2] = i[32];
  assign o[1] = i[16];
  assign o[0] = i[0];

endmodule

