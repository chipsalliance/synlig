module top;
   initial begin
      $display("Hex number ab should be printed: %h", 8'hAB);
   end
endmodule
