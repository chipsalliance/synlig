module top(output int o);
   int __FUNCTION__ = 15;
   assign o = __FUNCTION__;
endmodule
