

module top
(
  i,
  o
);

  input [1023:0] i;
  output [1023:0] o;

  bsg_array_reverse
  wrapper
  (
    .i(i),
    .o(o)
  );


endmodule



module bsg_array_reverse
(
  i,
  o
);

  input [1023:0] i;
  output [1023:0] o;
  wire [1023:0] o;
  assign o[1023] = i[15];
  assign o[1022] = i[14];
  assign o[1021] = i[13];
  assign o[1020] = i[12];
  assign o[1019] = i[11];
  assign o[1018] = i[10];
  assign o[1017] = i[9];
  assign o[1016] = i[8];
  assign o[1015] = i[7];
  assign o[1014] = i[6];
  assign o[1013] = i[5];
  assign o[1012] = i[4];
  assign o[1011] = i[3];
  assign o[1010] = i[2];
  assign o[1009] = i[1];
  assign o[1008] = i[0];
  assign o[1007] = i[31];
  assign o[1006] = i[30];
  assign o[1005] = i[29];
  assign o[1004] = i[28];
  assign o[1003] = i[27];
  assign o[1002] = i[26];
  assign o[1001] = i[25];
  assign o[1000] = i[24];
  assign o[999] = i[23];
  assign o[998] = i[22];
  assign o[997] = i[21];
  assign o[996] = i[20];
  assign o[995] = i[19];
  assign o[994] = i[18];
  assign o[993] = i[17];
  assign o[992] = i[16];
  assign o[991] = i[47];
  assign o[990] = i[46];
  assign o[989] = i[45];
  assign o[988] = i[44];
  assign o[987] = i[43];
  assign o[986] = i[42];
  assign o[985] = i[41];
  assign o[984] = i[40];
  assign o[983] = i[39];
  assign o[982] = i[38];
  assign o[981] = i[37];
  assign o[980] = i[36];
  assign o[979] = i[35];
  assign o[978] = i[34];
  assign o[977] = i[33];
  assign o[976] = i[32];
  assign o[975] = i[63];
  assign o[974] = i[62];
  assign o[973] = i[61];
  assign o[972] = i[60];
  assign o[971] = i[59];
  assign o[970] = i[58];
  assign o[969] = i[57];
  assign o[968] = i[56];
  assign o[967] = i[55];
  assign o[966] = i[54];
  assign o[965] = i[53];
  assign o[964] = i[52];
  assign o[963] = i[51];
  assign o[962] = i[50];
  assign o[961] = i[49];
  assign o[960] = i[48];
  assign o[959] = i[79];
  assign o[958] = i[78];
  assign o[957] = i[77];
  assign o[956] = i[76];
  assign o[955] = i[75];
  assign o[954] = i[74];
  assign o[953] = i[73];
  assign o[952] = i[72];
  assign o[951] = i[71];
  assign o[950] = i[70];
  assign o[949] = i[69];
  assign o[948] = i[68];
  assign o[947] = i[67];
  assign o[946] = i[66];
  assign o[945] = i[65];
  assign o[944] = i[64];
  assign o[943] = i[95];
  assign o[942] = i[94];
  assign o[941] = i[93];
  assign o[940] = i[92];
  assign o[939] = i[91];
  assign o[938] = i[90];
  assign o[937] = i[89];
  assign o[936] = i[88];
  assign o[935] = i[87];
  assign o[934] = i[86];
  assign o[933] = i[85];
  assign o[932] = i[84];
  assign o[931] = i[83];
  assign o[930] = i[82];
  assign o[929] = i[81];
  assign o[928] = i[80];
  assign o[927] = i[111];
  assign o[926] = i[110];
  assign o[925] = i[109];
  assign o[924] = i[108];
  assign o[923] = i[107];
  assign o[922] = i[106];
  assign o[921] = i[105];
  assign o[920] = i[104];
  assign o[919] = i[103];
  assign o[918] = i[102];
  assign o[917] = i[101];
  assign o[916] = i[100];
  assign o[915] = i[99];
  assign o[914] = i[98];
  assign o[913] = i[97];
  assign o[912] = i[96];
  assign o[911] = i[127];
  assign o[910] = i[126];
  assign o[909] = i[125];
  assign o[908] = i[124];
  assign o[907] = i[123];
  assign o[906] = i[122];
  assign o[905] = i[121];
  assign o[904] = i[120];
  assign o[903] = i[119];
  assign o[902] = i[118];
  assign o[901] = i[117];
  assign o[900] = i[116];
  assign o[899] = i[115];
  assign o[898] = i[114];
  assign o[897] = i[113];
  assign o[896] = i[112];
  assign o[895] = i[143];
  assign o[894] = i[142];
  assign o[893] = i[141];
  assign o[892] = i[140];
  assign o[891] = i[139];
  assign o[890] = i[138];
  assign o[889] = i[137];
  assign o[888] = i[136];
  assign o[887] = i[135];
  assign o[886] = i[134];
  assign o[885] = i[133];
  assign o[884] = i[132];
  assign o[883] = i[131];
  assign o[882] = i[130];
  assign o[881] = i[129];
  assign o[880] = i[128];
  assign o[879] = i[159];
  assign o[878] = i[158];
  assign o[877] = i[157];
  assign o[876] = i[156];
  assign o[875] = i[155];
  assign o[874] = i[154];
  assign o[873] = i[153];
  assign o[872] = i[152];
  assign o[871] = i[151];
  assign o[870] = i[150];
  assign o[869] = i[149];
  assign o[868] = i[148];
  assign o[867] = i[147];
  assign o[866] = i[146];
  assign o[865] = i[145];
  assign o[864] = i[144];
  assign o[863] = i[175];
  assign o[862] = i[174];
  assign o[861] = i[173];
  assign o[860] = i[172];
  assign o[859] = i[171];
  assign o[858] = i[170];
  assign o[857] = i[169];
  assign o[856] = i[168];
  assign o[855] = i[167];
  assign o[854] = i[166];
  assign o[853] = i[165];
  assign o[852] = i[164];
  assign o[851] = i[163];
  assign o[850] = i[162];
  assign o[849] = i[161];
  assign o[848] = i[160];
  assign o[847] = i[191];
  assign o[846] = i[190];
  assign o[845] = i[189];
  assign o[844] = i[188];
  assign o[843] = i[187];
  assign o[842] = i[186];
  assign o[841] = i[185];
  assign o[840] = i[184];
  assign o[839] = i[183];
  assign o[838] = i[182];
  assign o[837] = i[181];
  assign o[836] = i[180];
  assign o[835] = i[179];
  assign o[834] = i[178];
  assign o[833] = i[177];
  assign o[832] = i[176];
  assign o[831] = i[207];
  assign o[830] = i[206];
  assign o[829] = i[205];
  assign o[828] = i[204];
  assign o[827] = i[203];
  assign o[826] = i[202];
  assign o[825] = i[201];
  assign o[824] = i[200];
  assign o[823] = i[199];
  assign o[822] = i[198];
  assign o[821] = i[197];
  assign o[820] = i[196];
  assign o[819] = i[195];
  assign o[818] = i[194];
  assign o[817] = i[193];
  assign o[816] = i[192];
  assign o[815] = i[223];
  assign o[814] = i[222];
  assign o[813] = i[221];
  assign o[812] = i[220];
  assign o[811] = i[219];
  assign o[810] = i[218];
  assign o[809] = i[217];
  assign o[808] = i[216];
  assign o[807] = i[215];
  assign o[806] = i[214];
  assign o[805] = i[213];
  assign o[804] = i[212];
  assign o[803] = i[211];
  assign o[802] = i[210];
  assign o[801] = i[209];
  assign o[800] = i[208];
  assign o[799] = i[239];
  assign o[798] = i[238];
  assign o[797] = i[237];
  assign o[796] = i[236];
  assign o[795] = i[235];
  assign o[794] = i[234];
  assign o[793] = i[233];
  assign o[792] = i[232];
  assign o[791] = i[231];
  assign o[790] = i[230];
  assign o[789] = i[229];
  assign o[788] = i[228];
  assign o[787] = i[227];
  assign o[786] = i[226];
  assign o[785] = i[225];
  assign o[784] = i[224];
  assign o[783] = i[255];
  assign o[782] = i[254];
  assign o[781] = i[253];
  assign o[780] = i[252];
  assign o[779] = i[251];
  assign o[778] = i[250];
  assign o[777] = i[249];
  assign o[776] = i[248];
  assign o[775] = i[247];
  assign o[774] = i[246];
  assign o[773] = i[245];
  assign o[772] = i[244];
  assign o[771] = i[243];
  assign o[770] = i[242];
  assign o[769] = i[241];
  assign o[768] = i[240];
  assign o[767] = i[271];
  assign o[766] = i[270];
  assign o[765] = i[269];
  assign o[764] = i[268];
  assign o[763] = i[267];
  assign o[762] = i[266];
  assign o[761] = i[265];
  assign o[760] = i[264];
  assign o[759] = i[263];
  assign o[758] = i[262];
  assign o[757] = i[261];
  assign o[756] = i[260];
  assign o[755] = i[259];
  assign o[754] = i[258];
  assign o[753] = i[257];
  assign o[752] = i[256];
  assign o[751] = i[287];
  assign o[750] = i[286];
  assign o[749] = i[285];
  assign o[748] = i[284];
  assign o[747] = i[283];
  assign o[746] = i[282];
  assign o[745] = i[281];
  assign o[744] = i[280];
  assign o[743] = i[279];
  assign o[742] = i[278];
  assign o[741] = i[277];
  assign o[740] = i[276];
  assign o[739] = i[275];
  assign o[738] = i[274];
  assign o[737] = i[273];
  assign o[736] = i[272];
  assign o[735] = i[303];
  assign o[734] = i[302];
  assign o[733] = i[301];
  assign o[732] = i[300];
  assign o[731] = i[299];
  assign o[730] = i[298];
  assign o[729] = i[297];
  assign o[728] = i[296];
  assign o[727] = i[295];
  assign o[726] = i[294];
  assign o[725] = i[293];
  assign o[724] = i[292];
  assign o[723] = i[291];
  assign o[722] = i[290];
  assign o[721] = i[289];
  assign o[720] = i[288];
  assign o[719] = i[319];
  assign o[718] = i[318];
  assign o[717] = i[317];
  assign o[716] = i[316];
  assign o[715] = i[315];
  assign o[714] = i[314];
  assign o[713] = i[313];
  assign o[712] = i[312];
  assign o[711] = i[311];
  assign o[710] = i[310];
  assign o[709] = i[309];
  assign o[708] = i[308];
  assign o[707] = i[307];
  assign o[706] = i[306];
  assign o[705] = i[305];
  assign o[704] = i[304];
  assign o[703] = i[335];
  assign o[702] = i[334];
  assign o[701] = i[333];
  assign o[700] = i[332];
  assign o[699] = i[331];
  assign o[698] = i[330];
  assign o[697] = i[329];
  assign o[696] = i[328];
  assign o[695] = i[327];
  assign o[694] = i[326];
  assign o[693] = i[325];
  assign o[692] = i[324];
  assign o[691] = i[323];
  assign o[690] = i[322];
  assign o[689] = i[321];
  assign o[688] = i[320];
  assign o[687] = i[351];
  assign o[686] = i[350];
  assign o[685] = i[349];
  assign o[684] = i[348];
  assign o[683] = i[347];
  assign o[682] = i[346];
  assign o[681] = i[345];
  assign o[680] = i[344];
  assign o[679] = i[343];
  assign o[678] = i[342];
  assign o[677] = i[341];
  assign o[676] = i[340];
  assign o[675] = i[339];
  assign o[674] = i[338];
  assign o[673] = i[337];
  assign o[672] = i[336];
  assign o[671] = i[367];
  assign o[670] = i[366];
  assign o[669] = i[365];
  assign o[668] = i[364];
  assign o[667] = i[363];
  assign o[666] = i[362];
  assign o[665] = i[361];
  assign o[664] = i[360];
  assign o[663] = i[359];
  assign o[662] = i[358];
  assign o[661] = i[357];
  assign o[660] = i[356];
  assign o[659] = i[355];
  assign o[658] = i[354];
  assign o[657] = i[353];
  assign o[656] = i[352];
  assign o[655] = i[383];
  assign o[654] = i[382];
  assign o[653] = i[381];
  assign o[652] = i[380];
  assign o[651] = i[379];
  assign o[650] = i[378];
  assign o[649] = i[377];
  assign o[648] = i[376];
  assign o[647] = i[375];
  assign o[646] = i[374];
  assign o[645] = i[373];
  assign o[644] = i[372];
  assign o[643] = i[371];
  assign o[642] = i[370];
  assign o[641] = i[369];
  assign o[640] = i[368];
  assign o[639] = i[399];
  assign o[638] = i[398];
  assign o[637] = i[397];
  assign o[636] = i[396];
  assign o[635] = i[395];
  assign o[634] = i[394];
  assign o[633] = i[393];
  assign o[632] = i[392];
  assign o[631] = i[391];
  assign o[630] = i[390];
  assign o[629] = i[389];
  assign o[628] = i[388];
  assign o[627] = i[387];
  assign o[626] = i[386];
  assign o[625] = i[385];
  assign o[624] = i[384];
  assign o[623] = i[415];
  assign o[622] = i[414];
  assign o[621] = i[413];
  assign o[620] = i[412];
  assign o[619] = i[411];
  assign o[618] = i[410];
  assign o[617] = i[409];
  assign o[616] = i[408];
  assign o[615] = i[407];
  assign o[614] = i[406];
  assign o[613] = i[405];
  assign o[612] = i[404];
  assign o[611] = i[403];
  assign o[610] = i[402];
  assign o[609] = i[401];
  assign o[608] = i[400];
  assign o[607] = i[431];
  assign o[606] = i[430];
  assign o[605] = i[429];
  assign o[604] = i[428];
  assign o[603] = i[427];
  assign o[602] = i[426];
  assign o[601] = i[425];
  assign o[600] = i[424];
  assign o[599] = i[423];
  assign o[598] = i[422];
  assign o[597] = i[421];
  assign o[596] = i[420];
  assign o[595] = i[419];
  assign o[594] = i[418];
  assign o[593] = i[417];
  assign o[592] = i[416];
  assign o[591] = i[447];
  assign o[590] = i[446];
  assign o[589] = i[445];
  assign o[588] = i[444];
  assign o[587] = i[443];
  assign o[586] = i[442];
  assign o[585] = i[441];
  assign o[584] = i[440];
  assign o[583] = i[439];
  assign o[582] = i[438];
  assign o[581] = i[437];
  assign o[580] = i[436];
  assign o[579] = i[435];
  assign o[578] = i[434];
  assign o[577] = i[433];
  assign o[576] = i[432];
  assign o[575] = i[463];
  assign o[574] = i[462];
  assign o[573] = i[461];
  assign o[572] = i[460];
  assign o[571] = i[459];
  assign o[570] = i[458];
  assign o[569] = i[457];
  assign o[568] = i[456];
  assign o[567] = i[455];
  assign o[566] = i[454];
  assign o[565] = i[453];
  assign o[564] = i[452];
  assign o[563] = i[451];
  assign o[562] = i[450];
  assign o[561] = i[449];
  assign o[560] = i[448];
  assign o[559] = i[479];
  assign o[558] = i[478];
  assign o[557] = i[477];
  assign o[556] = i[476];
  assign o[555] = i[475];
  assign o[554] = i[474];
  assign o[553] = i[473];
  assign o[552] = i[472];
  assign o[551] = i[471];
  assign o[550] = i[470];
  assign o[549] = i[469];
  assign o[548] = i[468];
  assign o[547] = i[467];
  assign o[546] = i[466];
  assign o[545] = i[465];
  assign o[544] = i[464];
  assign o[543] = i[495];
  assign o[542] = i[494];
  assign o[541] = i[493];
  assign o[540] = i[492];
  assign o[539] = i[491];
  assign o[538] = i[490];
  assign o[537] = i[489];
  assign o[536] = i[488];
  assign o[535] = i[487];
  assign o[534] = i[486];
  assign o[533] = i[485];
  assign o[532] = i[484];
  assign o[531] = i[483];
  assign o[530] = i[482];
  assign o[529] = i[481];
  assign o[528] = i[480];
  assign o[527] = i[511];
  assign o[526] = i[510];
  assign o[525] = i[509];
  assign o[524] = i[508];
  assign o[523] = i[507];
  assign o[522] = i[506];
  assign o[521] = i[505];
  assign o[520] = i[504];
  assign o[519] = i[503];
  assign o[518] = i[502];
  assign o[517] = i[501];
  assign o[516] = i[500];
  assign o[515] = i[499];
  assign o[514] = i[498];
  assign o[513] = i[497];
  assign o[512] = i[496];
  assign o[511] = i[527];
  assign o[510] = i[526];
  assign o[509] = i[525];
  assign o[508] = i[524];
  assign o[507] = i[523];
  assign o[506] = i[522];
  assign o[505] = i[521];
  assign o[504] = i[520];
  assign o[503] = i[519];
  assign o[502] = i[518];
  assign o[501] = i[517];
  assign o[500] = i[516];
  assign o[499] = i[515];
  assign o[498] = i[514];
  assign o[497] = i[513];
  assign o[496] = i[512];
  assign o[495] = i[543];
  assign o[494] = i[542];
  assign o[493] = i[541];
  assign o[492] = i[540];
  assign o[491] = i[539];
  assign o[490] = i[538];
  assign o[489] = i[537];
  assign o[488] = i[536];
  assign o[487] = i[535];
  assign o[486] = i[534];
  assign o[485] = i[533];
  assign o[484] = i[532];
  assign o[483] = i[531];
  assign o[482] = i[530];
  assign o[481] = i[529];
  assign o[480] = i[528];
  assign o[479] = i[559];
  assign o[478] = i[558];
  assign o[477] = i[557];
  assign o[476] = i[556];
  assign o[475] = i[555];
  assign o[474] = i[554];
  assign o[473] = i[553];
  assign o[472] = i[552];
  assign o[471] = i[551];
  assign o[470] = i[550];
  assign o[469] = i[549];
  assign o[468] = i[548];
  assign o[467] = i[547];
  assign o[466] = i[546];
  assign o[465] = i[545];
  assign o[464] = i[544];
  assign o[463] = i[575];
  assign o[462] = i[574];
  assign o[461] = i[573];
  assign o[460] = i[572];
  assign o[459] = i[571];
  assign o[458] = i[570];
  assign o[457] = i[569];
  assign o[456] = i[568];
  assign o[455] = i[567];
  assign o[454] = i[566];
  assign o[453] = i[565];
  assign o[452] = i[564];
  assign o[451] = i[563];
  assign o[450] = i[562];
  assign o[449] = i[561];
  assign o[448] = i[560];
  assign o[447] = i[591];
  assign o[446] = i[590];
  assign o[445] = i[589];
  assign o[444] = i[588];
  assign o[443] = i[587];
  assign o[442] = i[586];
  assign o[441] = i[585];
  assign o[440] = i[584];
  assign o[439] = i[583];
  assign o[438] = i[582];
  assign o[437] = i[581];
  assign o[436] = i[580];
  assign o[435] = i[579];
  assign o[434] = i[578];
  assign o[433] = i[577];
  assign o[432] = i[576];
  assign o[431] = i[607];
  assign o[430] = i[606];
  assign o[429] = i[605];
  assign o[428] = i[604];
  assign o[427] = i[603];
  assign o[426] = i[602];
  assign o[425] = i[601];
  assign o[424] = i[600];
  assign o[423] = i[599];
  assign o[422] = i[598];
  assign o[421] = i[597];
  assign o[420] = i[596];
  assign o[419] = i[595];
  assign o[418] = i[594];
  assign o[417] = i[593];
  assign o[416] = i[592];
  assign o[415] = i[623];
  assign o[414] = i[622];
  assign o[413] = i[621];
  assign o[412] = i[620];
  assign o[411] = i[619];
  assign o[410] = i[618];
  assign o[409] = i[617];
  assign o[408] = i[616];
  assign o[407] = i[615];
  assign o[406] = i[614];
  assign o[405] = i[613];
  assign o[404] = i[612];
  assign o[403] = i[611];
  assign o[402] = i[610];
  assign o[401] = i[609];
  assign o[400] = i[608];
  assign o[399] = i[639];
  assign o[398] = i[638];
  assign o[397] = i[637];
  assign o[396] = i[636];
  assign o[395] = i[635];
  assign o[394] = i[634];
  assign o[393] = i[633];
  assign o[392] = i[632];
  assign o[391] = i[631];
  assign o[390] = i[630];
  assign o[389] = i[629];
  assign o[388] = i[628];
  assign o[387] = i[627];
  assign o[386] = i[626];
  assign o[385] = i[625];
  assign o[384] = i[624];
  assign o[383] = i[655];
  assign o[382] = i[654];
  assign o[381] = i[653];
  assign o[380] = i[652];
  assign o[379] = i[651];
  assign o[378] = i[650];
  assign o[377] = i[649];
  assign o[376] = i[648];
  assign o[375] = i[647];
  assign o[374] = i[646];
  assign o[373] = i[645];
  assign o[372] = i[644];
  assign o[371] = i[643];
  assign o[370] = i[642];
  assign o[369] = i[641];
  assign o[368] = i[640];
  assign o[367] = i[671];
  assign o[366] = i[670];
  assign o[365] = i[669];
  assign o[364] = i[668];
  assign o[363] = i[667];
  assign o[362] = i[666];
  assign o[361] = i[665];
  assign o[360] = i[664];
  assign o[359] = i[663];
  assign o[358] = i[662];
  assign o[357] = i[661];
  assign o[356] = i[660];
  assign o[355] = i[659];
  assign o[354] = i[658];
  assign o[353] = i[657];
  assign o[352] = i[656];
  assign o[351] = i[687];
  assign o[350] = i[686];
  assign o[349] = i[685];
  assign o[348] = i[684];
  assign o[347] = i[683];
  assign o[346] = i[682];
  assign o[345] = i[681];
  assign o[344] = i[680];
  assign o[343] = i[679];
  assign o[342] = i[678];
  assign o[341] = i[677];
  assign o[340] = i[676];
  assign o[339] = i[675];
  assign o[338] = i[674];
  assign o[337] = i[673];
  assign o[336] = i[672];
  assign o[335] = i[703];
  assign o[334] = i[702];
  assign o[333] = i[701];
  assign o[332] = i[700];
  assign o[331] = i[699];
  assign o[330] = i[698];
  assign o[329] = i[697];
  assign o[328] = i[696];
  assign o[327] = i[695];
  assign o[326] = i[694];
  assign o[325] = i[693];
  assign o[324] = i[692];
  assign o[323] = i[691];
  assign o[322] = i[690];
  assign o[321] = i[689];
  assign o[320] = i[688];
  assign o[319] = i[719];
  assign o[318] = i[718];
  assign o[317] = i[717];
  assign o[316] = i[716];
  assign o[315] = i[715];
  assign o[314] = i[714];
  assign o[313] = i[713];
  assign o[312] = i[712];
  assign o[311] = i[711];
  assign o[310] = i[710];
  assign o[309] = i[709];
  assign o[308] = i[708];
  assign o[307] = i[707];
  assign o[306] = i[706];
  assign o[305] = i[705];
  assign o[304] = i[704];
  assign o[303] = i[735];
  assign o[302] = i[734];
  assign o[301] = i[733];
  assign o[300] = i[732];
  assign o[299] = i[731];
  assign o[298] = i[730];
  assign o[297] = i[729];
  assign o[296] = i[728];
  assign o[295] = i[727];
  assign o[294] = i[726];
  assign o[293] = i[725];
  assign o[292] = i[724];
  assign o[291] = i[723];
  assign o[290] = i[722];
  assign o[289] = i[721];
  assign o[288] = i[720];
  assign o[287] = i[751];
  assign o[286] = i[750];
  assign o[285] = i[749];
  assign o[284] = i[748];
  assign o[283] = i[747];
  assign o[282] = i[746];
  assign o[281] = i[745];
  assign o[280] = i[744];
  assign o[279] = i[743];
  assign o[278] = i[742];
  assign o[277] = i[741];
  assign o[276] = i[740];
  assign o[275] = i[739];
  assign o[274] = i[738];
  assign o[273] = i[737];
  assign o[272] = i[736];
  assign o[271] = i[767];
  assign o[270] = i[766];
  assign o[269] = i[765];
  assign o[268] = i[764];
  assign o[267] = i[763];
  assign o[266] = i[762];
  assign o[265] = i[761];
  assign o[264] = i[760];
  assign o[263] = i[759];
  assign o[262] = i[758];
  assign o[261] = i[757];
  assign o[260] = i[756];
  assign o[259] = i[755];
  assign o[258] = i[754];
  assign o[257] = i[753];
  assign o[256] = i[752];
  assign o[255] = i[783];
  assign o[254] = i[782];
  assign o[253] = i[781];
  assign o[252] = i[780];
  assign o[251] = i[779];
  assign o[250] = i[778];
  assign o[249] = i[777];
  assign o[248] = i[776];
  assign o[247] = i[775];
  assign o[246] = i[774];
  assign o[245] = i[773];
  assign o[244] = i[772];
  assign o[243] = i[771];
  assign o[242] = i[770];
  assign o[241] = i[769];
  assign o[240] = i[768];
  assign o[239] = i[799];
  assign o[238] = i[798];
  assign o[237] = i[797];
  assign o[236] = i[796];
  assign o[235] = i[795];
  assign o[234] = i[794];
  assign o[233] = i[793];
  assign o[232] = i[792];
  assign o[231] = i[791];
  assign o[230] = i[790];
  assign o[229] = i[789];
  assign o[228] = i[788];
  assign o[227] = i[787];
  assign o[226] = i[786];
  assign o[225] = i[785];
  assign o[224] = i[784];
  assign o[223] = i[815];
  assign o[222] = i[814];
  assign o[221] = i[813];
  assign o[220] = i[812];
  assign o[219] = i[811];
  assign o[218] = i[810];
  assign o[217] = i[809];
  assign o[216] = i[808];
  assign o[215] = i[807];
  assign o[214] = i[806];
  assign o[213] = i[805];
  assign o[212] = i[804];
  assign o[211] = i[803];
  assign o[210] = i[802];
  assign o[209] = i[801];
  assign o[208] = i[800];
  assign o[207] = i[831];
  assign o[206] = i[830];
  assign o[205] = i[829];
  assign o[204] = i[828];
  assign o[203] = i[827];
  assign o[202] = i[826];
  assign o[201] = i[825];
  assign o[200] = i[824];
  assign o[199] = i[823];
  assign o[198] = i[822];
  assign o[197] = i[821];
  assign o[196] = i[820];
  assign o[195] = i[819];
  assign o[194] = i[818];
  assign o[193] = i[817];
  assign o[192] = i[816];
  assign o[191] = i[847];
  assign o[190] = i[846];
  assign o[189] = i[845];
  assign o[188] = i[844];
  assign o[187] = i[843];
  assign o[186] = i[842];
  assign o[185] = i[841];
  assign o[184] = i[840];
  assign o[183] = i[839];
  assign o[182] = i[838];
  assign o[181] = i[837];
  assign o[180] = i[836];
  assign o[179] = i[835];
  assign o[178] = i[834];
  assign o[177] = i[833];
  assign o[176] = i[832];
  assign o[175] = i[863];
  assign o[174] = i[862];
  assign o[173] = i[861];
  assign o[172] = i[860];
  assign o[171] = i[859];
  assign o[170] = i[858];
  assign o[169] = i[857];
  assign o[168] = i[856];
  assign o[167] = i[855];
  assign o[166] = i[854];
  assign o[165] = i[853];
  assign o[164] = i[852];
  assign o[163] = i[851];
  assign o[162] = i[850];
  assign o[161] = i[849];
  assign o[160] = i[848];
  assign o[159] = i[879];
  assign o[158] = i[878];
  assign o[157] = i[877];
  assign o[156] = i[876];
  assign o[155] = i[875];
  assign o[154] = i[874];
  assign o[153] = i[873];
  assign o[152] = i[872];
  assign o[151] = i[871];
  assign o[150] = i[870];
  assign o[149] = i[869];
  assign o[148] = i[868];
  assign o[147] = i[867];
  assign o[146] = i[866];
  assign o[145] = i[865];
  assign o[144] = i[864];
  assign o[143] = i[895];
  assign o[142] = i[894];
  assign o[141] = i[893];
  assign o[140] = i[892];
  assign o[139] = i[891];
  assign o[138] = i[890];
  assign o[137] = i[889];
  assign o[136] = i[888];
  assign o[135] = i[887];
  assign o[134] = i[886];
  assign o[133] = i[885];
  assign o[132] = i[884];
  assign o[131] = i[883];
  assign o[130] = i[882];
  assign o[129] = i[881];
  assign o[128] = i[880];
  assign o[127] = i[911];
  assign o[126] = i[910];
  assign o[125] = i[909];
  assign o[124] = i[908];
  assign o[123] = i[907];
  assign o[122] = i[906];
  assign o[121] = i[905];
  assign o[120] = i[904];
  assign o[119] = i[903];
  assign o[118] = i[902];
  assign o[117] = i[901];
  assign o[116] = i[900];
  assign o[115] = i[899];
  assign o[114] = i[898];
  assign o[113] = i[897];
  assign o[112] = i[896];
  assign o[111] = i[927];
  assign o[110] = i[926];
  assign o[109] = i[925];
  assign o[108] = i[924];
  assign o[107] = i[923];
  assign o[106] = i[922];
  assign o[105] = i[921];
  assign o[104] = i[920];
  assign o[103] = i[919];
  assign o[102] = i[918];
  assign o[101] = i[917];
  assign o[100] = i[916];
  assign o[99] = i[915];
  assign o[98] = i[914];
  assign o[97] = i[913];
  assign o[96] = i[912];
  assign o[95] = i[943];
  assign o[94] = i[942];
  assign o[93] = i[941];
  assign o[92] = i[940];
  assign o[91] = i[939];
  assign o[90] = i[938];
  assign o[89] = i[937];
  assign o[88] = i[936];
  assign o[87] = i[935];
  assign o[86] = i[934];
  assign o[85] = i[933];
  assign o[84] = i[932];
  assign o[83] = i[931];
  assign o[82] = i[930];
  assign o[81] = i[929];
  assign o[80] = i[928];
  assign o[79] = i[959];
  assign o[78] = i[958];
  assign o[77] = i[957];
  assign o[76] = i[956];
  assign o[75] = i[955];
  assign o[74] = i[954];
  assign o[73] = i[953];
  assign o[72] = i[952];
  assign o[71] = i[951];
  assign o[70] = i[950];
  assign o[69] = i[949];
  assign o[68] = i[948];
  assign o[67] = i[947];
  assign o[66] = i[946];
  assign o[65] = i[945];
  assign o[64] = i[944];
  assign o[63] = i[975];
  assign o[62] = i[974];
  assign o[61] = i[973];
  assign o[60] = i[972];
  assign o[59] = i[971];
  assign o[58] = i[970];
  assign o[57] = i[969];
  assign o[56] = i[968];
  assign o[55] = i[967];
  assign o[54] = i[966];
  assign o[53] = i[965];
  assign o[52] = i[964];
  assign o[51] = i[963];
  assign o[50] = i[962];
  assign o[49] = i[961];
  assign o[48] = i[960];
  assign o[47] = i[991];
  assign o[46] = i[990];
  assign o[45] = i[989];
  assign o[44] = i[988];
  assign o[43] = i[987];
  assign o[42] = i[986];
  assign o[41] = i[985];
  assign o[40] = i[984];
  assign o[39] = i[983];
  assign o[38] = i[982];
  assign o[37] = i[981];
  assign o[36] = i[980];
  assign o[35] = i[979];
  assign o[34] = i[978];
  assign o[33] = i[977];
  assign o[32] = i[976];
  assign o[31] = i[1007];
  assign o[30] = i[1006];
  assign o[29] = i[1005];
  assign o[28] = i[1004];
  assign o[27] = i[1003];
  assign o[26] = i[1002];
  assign o[25] = i[1001];
  assign o[24] = i[1000];
  assign o[23] = i[999];
  assign o[22] = i[998];
  assign o[21] = i[997];
  assign o[20] = i[996];
  assign o[19] = i[995];
  assign o[18] = i[994];
  assign o[17] = i[993];
  assign o[16] = i[992];
  assign o[15] = i[1023];
  assign o[14] = i[1022];
  assign o[13] = i[1021];
  assign o[12] = i[1020];
  assign o[11] = i[1019];
  assign o[10] = i[1018];
  assign o[9] = i[1017];
  assign o[8] = i[1016];
  assign o[7] = i[1015];
  assign o[6] = i[1014];
  assign o[5] = i[1013];
  assign o[4] = i[1012];
  assign o[3] = i[1011];
  assign o[2] = i[1010];
  assign o[1] = i[1009];
  assign o[0] = i[1008];

endmodule

