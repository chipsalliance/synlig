

module top
(
  clk_i,
  data_i,
  sel_i,
  data_o
);

  input [15:0] data_i;
  input [63:0] sel_i;
  output [15:0] data_o;
  input clk_i;

  bsg_fifo_shift_datapath
  wrapper
  (
    .data_i(data_i),
    .sel_i(sel_i),
    .data_o(data_o),
    .clk_i(clk_i)
  );


endmodule



module bsg_fifo_shift_datapath
(
  clk_i,
  data_i,
  sel_i,
  data_o
);

  input [15:0] data_i;
  input [63:0] sel_i;
  output [15:0] data_o;
  input clk_i;
  wire [15:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  r_31__15_,r_31__14_,r_31__13_,r_31__12_,r_31__11_,r_31__10_,r_31__9_,r_31__8_,
  r_31__7_,r_31__6_,r_31__5_,r_31__4_,r_31__3_,r_31__2_,r_31__1_,r_31__0_,r_30__15_,
  r_30__14_,r_30__13_,r_30__12_,r_30__11_,r_30__10_,r_30__9_,r_30__8_,r_30__7_,
  r_30__6_,r_30__5_,r_30__4_,r_30__3_,r_30__2_,r_30__1_,r_30__0_,r_29__15_,r_29__14_,
  r_29__13_,r_29__12_,r_29__11_,r_29__10_,r_29__9_,r_29__8_,r_29__7_,r_29__6_,
  r_29__5_,r_29__4_,r_29__3_,r_29__2_,r_29__1_,r_29__0_,r_28__15_,r_28__14_,r_28__13_,
  r_28__12_,r_28__11_,r_28__10_,r_28__9_,r_28__8_,r_28__7_,r_28__6_,r_28__5_,
  r_28__4_,r_28__3_,r_28__2_,r_28__1_,r_28__0_,r_27__15_,r_27__14_,r_27__13_,r_27__12_,
  r_27__11_,r_27__10_,r_27__9_,r_27__8_,r_27__7_,r_27__6_,r_27__5_,r_27__4_,
  r_27__3_,r_27__2_,r_27__1_,r_27__0_,r_26__15_,r_26__14_,r_26__13_,r_26__12_,r_26__11_,
  r_26__10_,r_26__9_,r_26__8_,r_26__7_,r_26__6_,r_26__5_,r_26__4_,r_26__3_,r_26__2_,
  r_26__1_,r_26__0_,r_25__15_,r_25__14_,r_25__13_,r_25__12_,r_25__11_,r_25__10_,
  r_25__9_,r_25__8_,r_25__7_,r_25__6_,r_25__5_,r_25__4_,r_25__3_,r_25__2_,r_25__1_,
  r_25__0_,r_24__15_,r_24__14_,r_24__13_,r_24__12_,r_24__11_,r_24__10_,r_24__9_,
  r_24__8_,r_24__7_,r_24__6_,r_24__5_,r_24__4_,r_24__3_,r_24__2_,r_24__1_,r_24__0_,
  r_23__15_,r_23__14_,r_23__13_,r_23__12_,r_23__11_,r_23__10_,r_23__9_,r_23__8_,
  r_23__7_,r_23__6_,r_23__5_,r_23__4_,r_23__3_,r_23__2_,r_23__1_,r_23__0_,r_22__15_,
  r_22__14_,r_22__13_,r_22__12_,r_22__11_,r_22__10_,r_22__9_,r_22__8_,r_22__7_,
  r_22__6_,r_22__5_,r_22__4_,r_22__3_,r_22__2_,r_22__1_,r_22__0_,r_21__15_,r_21__14_,
  r_21__13_,r_21__12_,r_21__11_,r_21__10_,r_21__9_,r_21__8_,r_21__7_,r_21__6_,
  r_21__5_,r_21__4_,r_21__3_,r_21__2_,r_21__1_,r_21__0_,r_20__15_,r_20__14_,r_20__13_,
  r_20__12_,r_20__11_,r_20__10_,r_20__9_,r_20__8_,r_20__7_,r_20__6_,r_20__5_,
  r_20__4_,r_20__3_,r_20__2_,r_20__1_,r_20__0_,r_19__15_,r_19__14_,r_19__13_,r_19__12_,
  r_19__11_,r_19__10_,r_19__9_,r_19__8_,r_19__7_,r_19__6_,r_19__5_,r_19__4_,
  r_19__3_,r_19__2_,r_19__1_,r_19__0_,r_18__15_,r_18__14_,r_18__13_,r_18__12_,r_18__11_,
  r_18__10_,r_18__9_,r_18__8_,r_18__7_,r_18__6_,r_18__5_,r_18__4_,r_18__3_,r_18__2_,
  r_18__1_,r_18__0_,r_17__15_,r_17__14_,r_17__13_,r_17__12_,r_17__11_,r_17__10_,
  r_17__9_,r_17__8_,r_17__7_,r_17__6_,r_17__5_,r_17__4_,r_17__3_,r_17__2_,r_17__1_,
  r_17__0_,r_16__15_,r_16__14_,r_16__13_,r_16__12_,r_16__11_,r_16__10_,r_16__9_,
  r_16__8_,r_16__7_,r_16__6_,r_16__5_,r_16__4_,r_16__3_,r_16__2_,r_16__1_,r_16__0_,
  r_15__15_,r_15__14_,r_15__13_,r_15__12_,r_15__11_,r_15__10_,r_15__9_,r_15__8_,
  r_15__7_,r_15__6_,r_15__5_,r_15__4_,r_15__3_,r_15__2_,r_15__1_,r_15__0_,r_14__15_,
  r_14__14_,r_14__13_,r_14__12_,r_14__11_,r_14__10_,r_14__9_,r_14__8_,r_14__7_,
  r_14__6_,r_14__5_,r_14__4_,r_14__3_,r_14__2_,r_14__1_,r_14__0_,r_13__15_,r_13__14_,
  r_13__13_,r_13__12_,r_13__11_,r_13__10_,r_13__9_,r_13__8_,r_13__7_,r_13__6_,
  r_13__5_,r_13__4_,r_13__3_,r_13__2_,r_13__1_,r_13__0_,r_12__15_,r_12__14_,r_12__13_,
  r_12__12_,r_12__11_,r_12__10_,r_12__9_,r_12__8_,r_12__7_,r_12__6_,r_12__5_,
  r_12__4_,r_12__3_,r_12__2_,r_12__1_,r_12__0_,r_11__15_,r_11__14_,r_11__13_,r_11__12_,
  r_11__11_,r_11__10_,r_11__9_,r_11__8_,r_11__7_,r_11__6_,r_11__5_,r_11__4_,
  r_11__3_,r_11__2_,r_11__1_,r_11__0_,r_10__15_,r_10__14_,r_10__13_,r_10__12_,r_10__11_,
  r_10__10_,r_10__9_,r_10__8_,r_10__7_,r_10__6_,r_10__5_,r_10__4_,r_10__3_,r_10__2_,
  r_10__1_,r_10__0_,r_9__15_,r_9__14_,r_9__13_,r_9__12_,r_9__11_,r_9__10_,r_9__9_,
  r_9__8_,r_9__7_,r_9__6_,r_9__5_,r_9__4_,r_9__3_,r_9__2_,r_9__1_,r_9__0_,
  r_8__15_,r_8__14_,r_8__13_,r_8__12_,r_8__11_,r_8__10_,r_8__9_,r_8__8_,r_8__7_,r_8__6_,
  r_8__5_,r_8__4_,r_8__3_,r_8__2_,r_8__1_,r_8__0_,r_7__15_,r_7__14_,r_7__13_,
  r_7__12_,r_7__11_,r_7__10_,r_7__9_,r_7__8_,r_7__7_,r_7__6_,r_7__5_,r_7__4_,r_7__3_,
  r_7__2_,r_7__1_,r_7__0_,r_6__15_,r_6__14_,r_6__13_,r_6__12_,r_6__11_,r_6__10_,
  r_6__9_,r_6__8_,r_6__7_,r_6__6_,r_6__5_,r_6__4_,r_6__3_,r_6__2_,r_6__1_,r_6__0_,
  r_5__15_,r_5__14_,r_5__13_,r_5__12_,r_5__11_,r_5__10_,r_5__9_,r_5__8_,r_5__7_,r_5__6_,
  r_5__5_,r_5__4_,r_5__3_,r_5__2_,r_5__1_,r_5__0_,r_4__15_,r_4__14_,r_4__13_,
  r_4__12_,r_4__11_,r_4__10_,r_4__9_,r_4__8_,r_4__7_,r_4__6_,r_4__5_,r_4__4_,r_4__3_,
  r_4__2_,r_4__1_,r_4__0_,r_3__15_,r_3__14_,r_3__13_,r_3__12_,r_3__11_,r_3__10_,
  r_3__9_,r_3__8_,r_3__7_,r_3__6_,r_3__5_,r_3__4_,r_3__3_,r_3__2_,r_3__1_,r_3__0_,
  r_2__15_,r_2__14_,r_2__13_,r_2__12_,r_2__11_,r_2__10_,r_2__9_,r_2__8_,r_2__7_,
  r_2__6_,r_2__5_,r_2__4_,r_2__3_,r_2__2_,r_2__1_,r_2__0_,r_1__15_,r_1__14_,r_1__13_,
  r_1__12_,r_1__11_,r_1__10_,r_1__9_,r_1__8_,r_1__7_,r_1__6_,r_1__5_,r_1__4_,r_1__3_,
  r_1__2_,r_1__1_,r_1__0_,N62,N63,N64,N65,N66,r_n_30__15_,r_n_30__14_,r_n_30__13_,
  r_n_30__12_,r_n_30__11_,r_n_30__10_,r_n_30__9_,r_n_30__8_,r_n_30__7_,r_n_30__6_,
  r_n_30__5_,r_n_30__4_,r_n_30__3_,r_n_30__2_,r_n_30__1_,r_n_30__0_,r_n_29__15_,
  r_n_29__14_,r_n_29__13_,r_n_29__12_,r_n_29__11_,r_n_29__10_,r_n_29__9_,r_n_29__8_,
  r_n_29__7_,r_n_29__6_,r_n_29__5_,r_n_29__4_,r_n_29__3_,r_n_29__2_,r_n_29__1_,
  r_n_29__0_,r_n_28__15_,r_n_28__14_,r_n_28__13_,r_n_28__12_,r_n_28__11_,r_n_28__10_,
  r_n_28__9_,r_n_28__8_,r_n_28__7_,r_n_28__6_,r_n_28__5_,r_n_28__4_,r_n_28__3_,
  r_n_28__2_,r_n_28__1_,r_n_28__0_,r_n_27__15_,r_n_27__14_,r_n_27__13_,r_n_27__12_,
  r_n_27__11_,r_n_27__10_,r_n_27__9_,r_n_27__8_,r_n_27__7_,r_n_27__6_,r_n_27__5_,
  r_n_27__4_,r_n_27__3_,r_n_27__2_,r_n_27__1_,r_n_27__0_,r_n_26__15_,r_n_26__14_,
  r_n_26__13_,r_n_26__12_,r_n_26__11_,r_n_26__10_,r_n_26__9_,r_n_26__8_,r_n_26__7_,
  r_n_26__6_,r_n_26__5_,r_n_26__4_,r_n_26__3_,r_n_26__2_,r_n_26__1_,r_n_26__0_,
  r_n_25__15_,r_n_25__14_,r_n_25__13_,r_n_25__12_,r_n_25__11_,r_n_25__10_,r_n_25__9_,
  r_n_25__8_,r_n_25__7_,r_n_25__6_,r_n_25__5_,r_n_25__4_,r_n_25__3_,r_n_25__2_,
  r_n_25__1_,r_n_25__0_,r_n_24__15_,r_n_24__14_,r_n_24__13_,r_n_24__12_,r_n_24__11_,
  r_n_24__10_,r_n_24__9_,r_n_24__8_,r_n_24__7_,r_n_24__6_,r_n_24__5_,r_n_24__4_,
  r_n_24__3_,r_n_24__2_,r_n_24__1_,r_n_24__0_,r_n_23__15_,r_n_23__14_,r_n_23__13_,
  r_n_23__12_,r_n_23__11_,r_n_23__10_,r_n_23__9_,r_n_23__8_,r_n_23__7_,r_n_23__6_,
  r_n_23__5_,r_n_23__4_,r_n_23__3_,r_n_23__2_,r_n_23__1_,r_n_23__0_,r_n_22__15_,
  r_n_22__14_,r_n_22__13_,r_n_22__12_,r_n_22__11_,r_n_22__10_,r_n_22__9_,r_n_22__8_,
  r_n_22__7_,r_n_22__6_,r_n_22__5_,r_n_22__4_,r_n_22__3_,r_n_22__2_,r_n_22__1_,
  r_n_22__0_,r_n_21__15_,r_n_21__14_,r_n_21__13_,r_n_21__12_,r_n_21__11_,r_n_21__10_,
  r_n_21__9_,r_n_21__8_,r_n_21__7_,r_n_21__6_,r_n_21__5_,r_n_21__4_,r_n_21__3_,
  r_n_21__2_,r_n_21__1_,r_n_21__0_,r_n_20__15_,r_n_20__14_,r_n_20__13_,r_n_20__12_,
  r_n_20__11_,r_n_20__10_,r_n_20__9_,r_n_20__8_,r_n_20__7_,r_n_20__6_,r_n_20__5_,
  r_n_20__4_,r_n_20__3_,r_n_20__2_,r_n_20__1_,r_n_20__0_,r_n_19__15_,r_n_19__14_,
  r_n_19__13_,r_n_19__12_,r_n_19__11_,r_n_19__10_,r_n_19__9_,r_n_19__8_,r_n_19__7_,
  r_n_19__6_,r_n_19__5_,r_n_19__4_,r_n_19__3_,r_n_19__2_,r_n_19__1_,r_n_19__0_,r_n_18__15_,
  r_n_18__14_,r_n_18__13_,r_n_18__12_,r_n_18__11_,r_n_18__10_,r_n_18__9_,
  r_n_18__8_,r_n_18__7_,r_n_18__6_,r_n_18__5_,r_n_18__4_,r_n_18__3_,r_n_18__2_,r_n_18__1_,
  r_n_18__0_,r_n_17__15_,r_n_17__14_,r_n_17__13_,r_n_17__12_,r_n_17__11_,
  r_n_17__10_,r_n_17__9_,r_n_17__8_,r_n_17__7_,r_n_17__6_,r_n_17__5_,r_n_17__4_,r_n_17__3_,
  r_n_17__2_,r_n_17__1_,r_n_17__0_,r_n_16__15_,r_n_16__14_,r_n_16__13_,r_n_16__12_,
  r_n_16__11_,r_n_16__10_,r_n_16__9_,r_n_16__8_,r_n_16__7_,r_n_16__6_,r_n_16__5_,
  r_n_16__4_,r_n_16__3_,r_n_16__2_,r_n_16__1_,r_n_16__0_,r_n_15__15_,r_n_15__14_,
  r_n_15__13_,r_n_15__12_,r_n_15__11_,r_n_15__10_,r_n_15__9_,r_n_15__8_,r_n_15__7_,
  r_n_15__6_,r_n_15__5_,r_n_15__4_,r_n_15__3_,r_n_15__2_,r_n_15__1_,r_n_15__0_,
  r_n_14__15_,r_n_14__14_,r_n_14__13_,r_n_14__12_,r_n_14__11_,r_n_14__10_,r_n_14__9_,
  r_n_14__8_,r_n_14__7_,r_n_14__6_,r_n_14__5_,r_n_14__4_,r_n_14__3_,r_n_14__2_,
  r_n_14__1_,r_n_14__0_,r_n_13__15_,r_n_13__14_,r_n_13__13_,r_n_13__12_,r_n_13__11_,
  r_n_13__10_,r_n_13__9_,r_n_13__8_,r_n_13__7_,r_n_13__6_,r_n_13__5_,r_n_13__4_,
  r_n_13__3_,r_n_13__2_,r_n_13__1_,r_n_13__0_,r_n_12__15_,r_n_12__14_,r_n_12__13_,
  r_n_12__12_,r_n_12__11_,r_n_12__10_,r_n_12__9_,r_n_12__8_,r_n_12__7_,r_n_12__6_,
  r_n_12__5_,r_n_12__4_,r_n_12__3_,r_n_12__2_,r_n_12__1_,r_n_12__0_,r_n_11__15_,
  r_n_11__14_,r_n_11__13_,r_n_11__12_,r_n_11__11_,r_n_11__10_,r_n_11__9_,r_n_11__8_,
  r_n_11__7_,r_n_11__6_,r_n_11__5_,r_n_11__4_,r_n_11__3_,r_n_11__2_,r_n_11__1_,
  r_n_11__0_,r_n_10__15_,r_n_10__14_,r_n_10__13_,r_n_10__12_,r_n_10__11_,r_n_10__10_,
  r_n_10__9_,r_n_10__8_,r_n_10__7_,r_n_10__6_,r_n_10__5_,r_n_10__4_,r_n_10__3_,
  r_n_10__2_,r_n_10__1_,r_n_10__0_,r_n_9__15_,r_n_9__14_,r_n_9__13_,r_n_9__12_,
  r_n_9__11_,r_n_9__10_,r_n_9__9_,r_n_9__8_,r_n_9__7_,r_n_9__6_,r_n_9__5_,r_n_9__4_,
  r_n_9__3_,r_n_9__2_,r_n_9__1_,r_n_9__0_,r_n_8__15_,r_n_8__14_,r_n_8__13_,r_n_8__12_,
  r_n_8__11_,r_n_8__10_,r_n_8__9_,r_n_8__8_,r_n_8__7_,r_n_8__6_,r_n_8__5_,r_n_8__4_,
  r_n_8__3_,r_n_8__2_,r_n_8__1_,r_n_8__0_,r_n_7__15_,r_n_7__14_,r_n_7__13_,
  r_n_7__12_,r_n_7__11_,r_n_7__10_,r_n_7__9_,r_n_7__8_,r_n_7__7_,r_n_7__6_,r_n_7__5_,
  r_n_7__4_,r_n_7__3_,r_n_7__2_,r_n_7__1_,r_n_7__0_,r_n_6__15_,r_n_6__14_,r_n_6__13_,
  r_n_6__12_,r_n_6__11_,r_n_6__10_,r_n_6__9_,r_n_6__8_,r_n_6__7_,r_n_6__6_,r_n_6__5_,
  r_n_6__4_,r_n_6__3_,r_n_6__2_,r_n_6__1_,r_n_6__0_,r_n_5__15_,r_n_5__14_,
  r_n_5__13_,r_n_5__12_,r_n_5__11_,r_n_5__10_,r_n_5__9_,r_n_5__8_,r_n_5__7_,r_n_5__6_,
  r_n_5__5_,r_n_5__4_,r_n_5__3_,r_n_5__2_,r_n_5__1_,r_n_5__0_,r_n_4__15_,r_n_4__14_,
  r_n_4__13_,r_n_4__12_,r_n_4__11_,r_n_4__10_,r_n_4__9_,r_n_4__8_,r_n_4__7_,
  r_n_4__6_,r_n_4__5_,r_n_4__4_,r_n_4__3_,r_n_4__2_,r_n_4__1_,r_n_4__0_,r_n_3__15_,
  r_n_3__14_,r_n_3__13_,r_n_3__12_,r_n_3__11_,r_n_3__10_,r_n_3__9_,r_n_3__8_,r_n_3__7_,
  r_n_3__6_,r_n_3__5_,r_n_3__4_,r_n_3__3_,r_n_3__2_,r_n_3__1_,r_n_3__0_,r_n_2__15_,
  r_n_2__14_,r_n_2__13_,r_n_2__12_,r_n_2__11_,r_n_2__10_,r_n_2__9_,r_n_2__8_,
  r_n_2__7_,r_n_2__6_,r_n_2__5_,r_n_2__4_,r_n_2__3_,r_n_2__2_,r_n_2__1_,r_n_2__0_,
  r_n_1__15_,r_n_1__14_,r_n_1__13_,r_n_1__12_,r_n_1__11_,r_n_1__10_,r_n_1__9_,r_n_1__8_,
  r_n_1__7_,r_n_1__6_,r_n_1__5_,r_n_1__4_,r_n_1__3_,r_n_1__2_,r_n_1__1_,r_n_1__0_,
  r_n_0__15_,r_n_0__14_,r_n_0__13_,r_n_0__12_,r_n_0__11_,r_n_0__10_,r_n_0__9_,
  r_n_0__8_,r_n_0__7_,r_n_0__6_,r_n_0__5_,r_n_0__4_,r_n_0__3_,r_n_0__2_,r_n_0__1_,
  r_n_0__0_,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,
  N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,
  N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,
  N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,
  N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,
  N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,
  N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,
  N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,
  N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,
  N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,
  N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,
  N248,N249,N250,N251,N252,N253,N254,N255;
  reg data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,
  data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,
  data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg,r_1__15__sv2v_reg,
  r_1__14__sv2v_reg,r_1__13__sv2v_reg,r_1__12__sv2v_reg,r_1__11__sv2v_reg,
  r_1__10__sv2v_reg,r_1__9__sv2v_reg,r_1__8__sv2v_reg,r_1__7__sv2v_reg,r_1__6__sv2v_reg,
  r_1__5__sv2v_reg,r_1__4__sv2v_reg,r_1__3__sv2v_reg,r_1__2__sv2v_reg,r_1__1__sv2v_reg,
  r_1__0__sv2v_reg,r_2__15__sv2v_reg,r_2__14__sv2v_reg,r_2__13__sv2v_reg,
  r_2__12__sv2v_reg,r_2__11__sv2v_reg,r_2__10__sv2v_reg,r_2__9__sv2v_reg,r_2__8__sv2v_reg,
  r_2__7__sv2v_reg,r_2__6__sv2v_reg,r_2__5__sv2v_reg,r_2__4__sv2v_reg,r_2__3__sv2v_reg,
  r_2__2__sv2v_reg,r_2__1__sv2v_reg,r_2__0__sv2v_reg,r_3__15__sv2v_reg,
  r_3__14__sv2v_reg,r_3__13__sv2v_reg,r_3__12__sv2v_reg,r_3__11__sv2v_reg,r_3__10__sv2v_reg,
  r_3__9__sv2v_reg,r_3__8__sv2v_reg,r_3__7__sv2v_reg,r_3__6__sv2v_reg,
  r_3__5__sv2v_reg,r_3__4__sv2v_reg,r_3__3__sv2v_reg,r_3__2__sv2v_reg,r_3__1__sv2v_reg,
  r_3__0__sv2v_reg,r_4__15__sv2v_reg,r_4__14__sv2v_reg,r_4__13__sv2v_reg,r_4__12__sv2v_reg,
  r_4__11__sv2v_reg,r_4__10__sv2v_reg,r_4__9__sv2v_reg,r_4__8__sv2v_reg,
  r_4__7__sv2v_reg,r_4__6__sv2v_reg,r_4__5__sv2v_reg,r_4__4__sv2v_reg,r_4__3__sv2v_reg,
  r_4__2__sv2v_reg,r_4__1__sv2v_reg,r_4__0__sv2v_reg,r_5__15__sv2v_reg,
  r_5__14__sv2v_reg,r_5__13__sv2v_reg,r_5__12__sv2v_reg,r_5__11__sv2v_reg,r_5__10__sv2v_reg,
  r_5__9__sv2v_reg,r_5__8__sv2v_reg,r_5__7__sv2v_reg,r_5__6__sv2v_reg,r_5__5__sv2v_reg,
  r_5__4__sv2v_reg,r_5__3__sv2v_reg,r_5__2__sv2v_reg,r_5__1__sv2v_reg,
  r_5__0__sv2v_reg,r_6__15__sv2v_reg,r_6__14__sv2v_reg,r_6__13__sv2v_reg,r_6__12__sv2v_reg,
  r_6__11__sv2v_reg,r_6__10__sv2v_reg,r_6__9__sv2v_reg,r_6__8__sv2v_reg,
  r_6__7__sv2v_reg,r_6__6__sv2v_reg,r_6__5__sv2v_reg,r_6__4__sv2v_reg,r_6__3__sv2v_reg,
  r_6__2__sv2v_reg,r_6__1__sv2v_reg,r_6__0__sv2v_reg,r_7__15__sv2v_reg,r_7__14__sv2v_reg,
  r_7__13__sv2v_reg,r_7__12__sv2v_reg,r_7__11__sv2v_reg,r_7__10__sv2v_reg,
  r_7__9__sv2v_reg,r_7__8__sv2v_reg,r_7__7__sv2v_reg,r_7__6__sv2v_reg,r_7__5__sv2v_reg,
  r_7__4__sv2v_reg,r_7__3__sv2v_reg,r_7__2__sv2v_reg,r_7__1__sv2v_reg,r_7__0__sv2v_reg,
  r_8__15__sv2v_reg,r_8__14__sv2v_reg,r_8__13__sv2v_reg,r_8__12__sv2v_reg,
  r_8__11__sv2v_reg,r_8__10__sv2v_reg,r_8__9__sv2v_reg,r_8__8__sv2v_reg,r_8__7__sv2v_reg,
  r_8__6__sv2v_reg,r_8__5__sv2v_reg,r_8__4__sv2v_reg,r_8__3__sv2v_reg,
  r_8__2__sv2v_reg,r_8__1__sv2v_reg,r_8__0__sv2v_reg,r_9__15__sv2v_reg,r_9__14__sv2v_reg,
  r_9__13__sv2v_reg,r_9__12__sv2v_reg,r_9__11__sv2v_reg,r_9__10__sv2v_reg,
  r_9__9__sv2v_reg,r_9__8__sv2v_reg,r_9__7__sv2v_reg,r_9__6__sv2v_reg,r_9__5__sv2v_reg,
  r_9__4__sv2v_reg,r_9__3__sv2v_reg,r_9__2__sv2v_reg,r_9__1__sv2v_reg,r_9__0__sv2v_reg,
  r_10__15__sv2v_reg,r_10__14__sv2v_reg,r_10__13__sv2v_reg,r_10__12__sv2v_reg,
  r_10__11__sv2v_reg,r_10__10__sv2v_reg,r_10__9__sv2v_reg,r_10__8__sv2v_reg,
  r_10__7__sv2v_reg,r_10__6__sv2v_reg,r_10__5__sv2v_reg,r_10__4__sv2v_reg,r_10__3__sv2v_reg,
  r_10__2__sv2v_reg,r_10__1__sv2v_reg,r_10__0__sv2v_reg,r_11__15__sv2v_reg,
  r_11__14__sv2v_reg,r_11__13__sv2v_reg,r_11__12__sv2v_reg,r_11__11__sv2v_reg,
  r_11__10__sv2v_reg,r_11__9__sv2v_reg,r_11__8__sv2v_reg,r_11__7__sv2v_reg,r_11__6__sv2v_reg,
  r_11__5__sv2v_reg,r_11__4__sv2v_reg,r_11__3__sv2v_reg,r_11__2__sv2v_reg,
  r_11__1__sv2v_reg,r_11__0__sv2v_reg,r_12__15__sv2v_reg,r_12__14__sv2v_reg,
  r_12__13__sv2v_reg,r_12__12__sv2v_reg,r_12__11__sv2v_reg,r_12__10__sv2v_reg,r_12__9__sv2v_reg,
  r_12__8__sv2v_reg,r_12__7__sv2v_reg,r_12__6__sv2v_reg,r_12__5__sv2v_reg,
  r_12__4__sv2v_reg,r_12__3__sv2v_reg,r_12__2__sv2v_reg,r_12__1__sv2v_reg,r_12__0__sv2v_reg,
  r_13__15__sv2v_reg,r_13__14__sv2v_reg,r_13__13__sv2v_reg,r_13__12__sv2v_reg,
  r_13__11__sv2v_reg,r_13__10__sv2v_reg,r_13__9__sv2v_reg,r_13__8__sv2v_reg,
  r_13__7__sv2v_reg,r_13__6__sv2v_reg,r_13__5__sv2v_reg,r_13__4__sv2v_reg,r_13__3__sv2v_reg,
  r_13__2__sv2v_reg,r_13__1__sv2v_reg,r_13__0__sv2v_reg,r_14__15__sv2v_reg,
  r_14__14__sv2v_reg,r_14__13__sv2v_reg,r_14__12__sv2v_reg,r_14__11__sv2v_reg,
  r_14__10__sv2v_reg,r_14__9__sv2v_reg,r_14__8__sv2v_reg,r_14__7__sv2v_reg,r_14__6__sv2v_reg,
  r_14__5__sv2v_reg,r_14__4__sv2v_reg,r_14__3__sv2v_reg,r_14__2__sv2v_reg,
  r_14__1__sv2v_reg,r_14__0__sv2v_reg,r_15__15__sv2v_reg,r_15__14__sv2v_reg,
  r_15__13__sv2v_reg,r_15__12__sv2v_reg,r_15__11__sv2v_reg,r_15__10__sv2v_reg,r_15__9__sv2v_reg,
  r_15__8__sv2v_reg,r_15__7__sv2v_reg,r_15__6__sv2v_reg,r_15__5__sv2v_reg,
  r_15__4__sv2v_reg,r_15__3__sv2v_reg,r_15__2__sv2v_reg,r_15__1__sv2v_reg,r_15__0__sv2v_reg,
  r_16__15__sv2v_reg,r_16__14__sv2v_reg,r_16__13__sv2v_reg,r_16__12__sv2v_reg,
  r_16__11__sv2v_reg,r_16__10__sv2v_reg,r_16__9__sv2v_reg,r_16__8__sv2v_reg,
  r_16__7__sv2v_reg,r_16__6__sv2v_reg,r_16__5__sv2v_reg,r_16__4__sv2v_reg,r_16__3__sv2v_reg,
  r_16__2__sv2v_reg,r_16__1__sv2v_reg,r_16__0__sv2v_reg,r_17__15__sv2v_reg,
  r_17__14__sv2v_reg,r_17__13__sv2v_reg,r_17__12__sv2v_reg,r_17__11__sv2v_reg,
  r_17__10__sv2v_reg,r_17__9__sv2v_reg,r_17__8__sv2v_reg,r_17__7__sv2v_reg,r_17__6__sv2v_reg,
  r_17__5__sv2v_reg,r_17__4__sv2v_reg,r_17__3__sv2v_reg,r_17__2__sv2v_reg,
  r_17__1__sv2v_reg,r_17__0__sv2v_reg,r_18__15__sv2v_reg,r_18__14__sv2v_reg,
  r_18__13__sv2v_reg,r_18__12__sv2v_reg,r_18__11__sv2v_reg,r_18__10__sv2v_reg,r_18__9__sv2v_reg,
  r_18__8__sv2v_reg,r_18__7__sv2v_reg,r_18__6__sv2v_reg,r_18__5__sv2v_reg,
  r_18__4__sv2v_reg,r_18__3__sv2v_reg,r_18__2__sv2v_reg,r_18__1__sv2v_reg,
  r_18__0__sv2v_reg,r_19__15__sv2v_reg,r_19__14__sv2v_reg,r_19__13__sv2v_reg,r_19__12__sv2v_reg,
  r_19__11__sv2v_reg,r_19__10__sv2v_reg,r_19__9__sv2v_reg,r_19__8__sv2v_reg,
  r_19__7__sv2v_reg,r_19__6__sv2v_reg,r_19__5__sv2v_reg,r_19__4__sv2v_reg,
  r_19__3__sv2v_reg,r_19__2__sv2v_reg,r_19__1__sv2v_reg,r_19__0__sv2v_reg,r_20__15__sv2v_reg,
  r_20__14__sv2v_reg,r_20__13__sv2v_reg,r_20__12__sv2v_reg,r_20__11__sv2v_reg,
  r_20__10__sv2v_reg,r_20__9__sv2v_reg,r_20__8__sv2v_reg,r_20__7__sv2v_reg,
  r_20__6__sv2v_reg,r_20__5__sv2v_reg,r_20__4__sv2v_reg,r_20__3__sv2v_reg,r_20__2__sv2v_reg,
  r_20__1__sv2v_reg,r_20__0__sv2v_reg,r_21__15__sv2v_reg,r_21__14__sv2v_reg,
  r_21__13__sv2v_reg,r_21__12__sv2v_reg,r_21__11__sv2v_reg,r_21__10__sv2v_reg,
  r_21__9__sv2v_reg,r_21__8__sv2v_reg,r_21__7__sv2v_reg,r_21__6__sv2v_reg,r_21__5__sv2v_reg,
  r_21__4__sv2v_reg,r_21__3__sv2v_reg,r_21__2__sv2v_reg,r_21__1__sv2v_reg,
  r_21__0__sv2v_reg,r_22__15__sv2v_reg,r_22__14__sv2v_reg,r_22__13__sv2v_reg,r_22__12__sv2v_reg,
  r_22__11__sv2v_reg,r_22__10__sv2v_reg,r_22__9__sv2v_reg,r_22__8__sv2v_reg,
  r_22__7__sv2v_reg,r_22__6__sv2v_reg,r_22__5__sv2v_reg,r_22__4__sv2v_reg,
  r_22__3__sv2v_reg,r_22__2__sv2v_reg,r_22__1__sv2v_reg,r_22__0__sv2v_reg,r_23__15__sv2v_reg,
  r_23__14__sv2v_reg,r_23__13__sv2v_reg,r_23__12__sv2v_reg,r_23__11__sv2v_reg,
  r_23__10__sv2v_reg,r_23__9__sv2v_reg,r_23__8__sv2v_reg,r_23__7__sv2v_reg,
  r_23__6__sv2v_reg,r_23__5__sv2v_reg,r_23__4__sv2v_reg,r_23__3__sv2v_reg,r_23__2__sv2v_reg,
  r_23__1__sv2v_reg,r_23__0__sv2v_reg,r_24__15__sv2v_reg,r_24__14__sv2v_reg,
  r_24__13__sv2v_reg,r_24__12__sv2v_reg,r_24__11__sv2v_reg,r_24__10__sv2v_reg,
  r_24__9__sv2v_reg,r_24__8__sv2v_reg,r_24__7__sv2v_reg,r_24__6__sv2v_reg,r_24__5__sv2v_reg,
  r_24__4__sv2v_reg,r_24__3__sv2v_reg,r_24__2__sv2v_reg,r_24__1__sv2v_reg,
  r_24__0__sv2v_reg,r_25__15__sv2v_reg,r_25__14__sv2v_reg,r_25__13__sv2v_reg,
  r_25__12__sv2v_reg,r_25__11__sv2v_reg,r_25__10__sv2v_reg,r_25__9__sv2v_reg,r_25__8__sv2v_reg,
  r_25__7__sv2v_reg,r_25__6__sv2v_reg,r_25__5__sv2v_reg,r_25__4__sv2v_reg,
  r_25__3__sv2v_reg,r_25__2__sv2v_reg,r_25__1__sv2v_reg,r_25__0__sv2v_reg,r_26__15__sv2v_reg,
  r_26__14__sv2v_reg,r_26__13__sv2v_reg,r_26__12__sv2v_reg,r_26__11__sv2v_reg,
  r_26__10__sv2v_reg,r_26__9__sv2v_reg,r_26__8__sv2v_reg,r_26__7__sv2v_reg,
  r_26__6__sv2v_reg,r_26__5__sv2v_reg,r_26__4__sv2v_reg,r_26__3__sv2v_reg,r_26__2__sv2v_reg,
  r_26__1__sv2v_reg,r_26__0__sv2v_reg,r_27__15__sv2v_reg,r_27__14__sv2v_reg,
  r_27__13__sv2v_reg,r_27__12__sv2v_reg,r_27__11__sv2v_reg,r_27__10__sv2v_reg,
  r_27__9__sv2v_reg,r_27__8__sv2v_reg,r_27__7__sv2v_reg,r_27__6__sv2v_reg,r_27__5__sv2v_reg,
  r_27__4__sv2v_reg,r_27__3__sv2v_reg,r_27__2__sv2v_reg,r_27__1__sv2v_reg,
  r_27__0__sv2v_reg,r_28__15__sv2v_reg,r_28__14__sv2v_reg,r_28__13__sv2v_reg,
  r_28__12__sv2v_reg,r_28__11__sv2v_reg,r_28__10__sv2v_reg,r_28__9__sv2v_reg,r_28__8__sv2v_reg,
  r_28__7__sv2v_reg,r_28__6__sv2v_reg,r_28__5__sv2v_reg,r_28__4__sv2v_reg,
  r_28__3__sv2v_reg,r_28__2__sv2v_reg,r_28__1__sv2v_reg,r_28__0__sv2v_reg,
  r_29__15__sv2v_reg,r_29__14__sv2v_reg,r_29__13__sv2v_reg,r_29__12__sv2v_reg,r_29__11__sv2v_reg,
  r_29__10__sv2v_reg,r_29__9__sv2v_reg,r_29__8__sv2v_reg,r_29__7__sv2v_reg,
  r_29__6__sv2v_reg,r_29__5__sv2v_reg,r_29__4__sv2v_reg,r_29__3__sv2v_reg,r_29__2__sv2v_reg,
  r_29__1__sv2v_reg,r_29__0__sv2v_reg,r_30__15__sv2v_reg,r_30__14__sv2v_reg,
  r_30__13__sv2v_reg,r_30__12__sv2v_reg,r_30__11__sv2v_reg,r_30__10__sv2v_reg,
  r_30__9__sv2v_reg,r_30__8__sv2v_reg,r_30__7__sv2v_reg,r_30__6__sv2v_reg,r_30__5__sv2v_reg,
  r_30__4__sv2v_reg,r_30__3__sv2v_reg,r_30__2__sv2v_reg,r_30__1__sv2v_reg,
  r_30__0__sv2v_reg,r_31__15__sv2v_reg,r_31__14__sv2v_reg,r_31__13__sv2v_reg,
  r_31__12__sv2v_reg,r_31__11__sv2v_reg,r_31__10__sv2v_reg,r_31__9__sv2v_reg,r_31__8__sv2v_reg,
  r_31__7__sv2v_reg,r_31__6__sv2v_reg,r_31__5__sv2v_reg,r_31__4__sv2v_reg,
  r_31__3__sv2v_reg,r_31__2__sv2v_reg,r_31__1__sv2v_reg,r_31__0__sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign r_1__15_ = r_1__15__sv2v_reg;
  assign r_1__14_ = r_1__14__sv2v_reg;
  assign r_1__13_ = r_1__13__sv2v_reg;
  assign r_1__12_ = r_1__12__sv2v_reg;
  assign r_1__11_ = r_1__11__sv2v_reg;
  assign r_1__10_ = r_1__10__sv2v_reg;
  assign r_1__9_ = r_1__9__sv2v_reg;
  assign r_1__8_ = r_1__8__sv2v_reg;
  assign r_1__7_ = r_1__7__sv2v_reg;
  assign r_1__6_ = r_1__6__sv2v_reg;
  assign r_1__5_ = r_1__5__sv2v_reg;
  assign r_1__4_ = r_1__4__sv2v_reg;
  assign r_1__3_ = r_1__3__sv2v_reg;
  assign r_1__2_ = r_1__2__sv2v_reg;
  assign r_1__1_ = r_1__1__sv2v_reg;
  assign r_1__0_ = r_1__0__sv2v_reg;
  assign r_2__15_ = r_2__15__sv2v_reg;
  assign r_2__14_ = r_2__14__sv2v_reg;
  assign r_2__13_ = r_2__13__sv2v_reg;
  assign r_2__12_ = r_2__12__sv2v_reg;
  assign r_2__11_ = r_2__11__sv2v_reg;
  assign r_2__10_ = r_2__10__sv2v_reg;
  assign r_2__9_ = r_2__9__sv2v_reg;
  assign r_2__8_ = r_2__8__sv2v_reg;
  assign r_2__7_ = r_2__7__sv2v_reg;
  assign r_2__6_ = r_2__6__sv2v_reg;
  assign r_2__5_ = r_2__5__sv2v_reg;
  assign r_2__4_ = r_2__4__sv2v_reg;
  assign r_2__3_ = r_2__3__sv2v_reg;
  assign r_2__2_ = r_2__2__sv2v_reg;
  assign r_2__1_ = r_2__1__sv2v_reg;
  assign r_2__0_ = r_2__0__sv2v_reg;
  assign r_3__15_ = r_3__15__sv2v_reg;
  assign r_3__14_ = r_3__14__sv2v_reg;
  assign r_3__13_ = r_3__13__sv2v_reg;
  assign r_3__12_ = r_3__12__sv2v_reg;
  assign r_3__11_ = r_3__11__sv2v_reg;
  assign r_3__10_ = r_3__10__sv2v_reg;
  assign r_3__9_ = r_3__9__sv2v_reg;
  assign r_3__8_ = r_3__8__sv2v_reg;
  assign r_3__7_ = r_3__7__sv2v_reg;
  assign r_3__6_ = r_3__6__sv2v_reg;
  assign r_3__5_ = r_3__5__sv2v_reg;
  assign r_3__4_ = r_3__4__sv2v_reg;
  assign r_3__3_ = r_3__3__sv2v_reg;
  assign r_3__2_ = r_3__2__sv2v_reg;
  assign r_3__1_ = r_3__1__sv2v_reg;
  assign r_3__0_ = r_3__0__sv2v_reg;
  assign r_4__15_ = r_4__15__sv2v_reg;
  assign r_4__14_ = r_4__14__sv2v_reg;
  assign r_4__13_ = r_4__13__sv2v_reg;
  assign r_4__12_ = r_4__12__sv2v_reg;
  assign r_4__11_ = r_4__11__sv2v_reg;
  assign r_4__10_ = r_4__10__sv2v_reg;
  assign r_4__9_ = r_4__9__sv2v_reg;
  assign r_4__8_ = r_4__8__sv2v_reg;
  assign r_4__7_ = r_4__7__sv2v_reg;
  assign r_4__6_ = r_4__6__sv2v_reg;
  assign r_4__5_ = r_4__5__sv2v_reg;
  assign r_4__4_ = r_4__4__sv2v_reg;
  assign r_4__3_ = r_4__3__sv2v_reg;
  assign r_4__2_ = r_4__2__sv2v_reg;
  assign r_4__1_ = r_4__1__sv2v_reg;
  assign r_4__0_ = r_4__0__sv2v_reg;
  assign r_5__15_ = r_5__15__sv2v_reg;
  assign r_5__14_ = r_5__14__sv2v_reg;
  assign r_5__13_ = r_5__13__sv2v_reg;
  assign r_5__12_ = r_5__12__sv2v_reg;
  assign r_5__11_ = r_5__11__sv2v_reg;
  assign r_5__10_ = r_5__10__sv2v_reg;
  assign r_5__9_ = r_5__9__sv2v_reg;
  assign r_5__8_ = r_5__8__sv2v_reg;
  assign r_5__7_ = r_5__7__sv2v_reg;
  assign r_5__6_ = r_5__6__sv2v_reg;
  assign r_5__5_ = r_5__5__sv2v_reg;
  assign r_5__4_ = r_5__4__sv2v_reg;
  assign r_5__3_ = r_5__3__sv2v_reg;
  assign r_5__2_ = r_5__2__sv2v_reg;
  assign r_5__1_ = r_5__1__sv2v_reg;
  assign r_5__0_ = r_5__0__sv2v_reg;
  assign r_6__15_ = r_6__15__sv2v_reg;
  assign r_6__14_ = r_6__14__sv2v_reg;
  assign r_6__13_ = r_6__13__sv2v_reg;
  assign r_6__12_ = r_6__12__sv2v_reg;
  assign r_6__11_ = r_6__11__sv2v_reg;
  assign r_6__10_ = r_6__10__sv2v_reg;
  assign r_6__9_ = r_6__9__sv2v_reg;
  assign r_6__8_ = r_6__8__sv2v_reg;
  assign r_6__7_ = r_6__7__sv2v_reg;
  assign r_6__6_ = r_6__6__sv2v_reg;
  assign r_6__5_ = r_6__5__sv2v_reg;
  assign r_6__4_ = r_6__4__sv2v_reg;
  assign r_6__3_ = r_6__3__sv2v_reg;
  assign r_6__2_ = r_6__2__sv2v_reg;
  assign r_6__1_ = r_6__1__sv2v_reg;
  assign r_6__0_ = r_6__0__sv2v_reg;
  assign r_7__15_ = r_7__15__sv2v_reg;
  assign r_7__14_ = r_7__14__sv2v_reg;
  assign r_7__13_ = r_7__13__sv2v_reg;
  assign r_7__12_ = r_7__12__sv2v_reg;
  assign r_7__11_ = r_7__11__sv2v_reg;
  assign r_7__10_ = r_7__10__sv2v_reg;
  assign r_7__9_ = r_7__9__sv2v_reg;
  assign r_7__8_ = r_7__8__sv2v_reg;
  assign r_7__7_ = r_7__7__sv2v_reg;
  assign r_7__6_ = r_7__6__sv2v_reg;
  assign r_7__5_ = r_7__5__sv2v_reg;
  assign r_7__4_ = r_7__4__sv2v_reg;
  assign r_7__3_ = r_7__3__sv2v_reg;
  assign r_7__2_ = r_7__2__sv2v_reg;
  assign r_7__1_ = r_7__1__sv2v_reg;
  assign r_7__0_ = r_7__0__sv2v_reg;
  assign r_8__15_ = r_8__15__sv2v_reg;
  assign r_8__14_ = r_8__14__sv2v_reg;
  assign r_8__13_ = r_8__13__sv2v_reg;
  assign r_8__12_ = r_8__12__sv2v_reg;
  assign r_8__11_ = r_8__11__sv2v_reg;
  assign r_8__10_ = r_8__10__sv2v_reg;
  assign r_8__9_ = r_8__9__sv2v_reg;
  assign r_8__8_ = r_8__8__sv2v_reg;
  assign r_8__7_ = r_8__7__sv2v_reg;
  assign r_8__6_ = r_8__6__sv2v_reg;
  assign r_8__5_ = r_8__5__sv2v_reg;
  assign r_8__4_ = r_8__4__sv2v_reg;
  assign r_8__3_ = r_8__3__sv2v_reg;
  assign r_8__2_ = r_8__2__sv2v_reg;
  assign r_8__1_ = r_8__1__sv2v_reg;
  assign r_8__0_ = r_8__0__sv2v_reg;
  assign r_9__15_ = r_9__15__sv2v_reg;
  assign r_9__14_ = r_9__14__sv2v_reg;
  assign r_9__13_ = r_9__13__sv2v_reg;
  assign r_9__12_ = r_9__12__sv2v_reg;
  assign r_9__11_ = r_9__11__sv2v_reg;
  assign r_9__10_ = r_9__10__sv2v_reg;
  assign r_9__9_ = r_9__9__sv2v_reg;
  assign r_9__8_ = r_9__8__sv2v_reg;
  assign r_9__7_ = r_9__7__sv2v_reg;
  assign r_9__6_ = r_9__6__sv2v_reg;
  assign r_9__5_ = r_9__5__sv2v_reg;
  assign r_9__4_ = r_9__4__sv2v_reg;
  assign r_9__3_ = r_9__3__sv2v_reg;
  assign r_9__2_ = r_9__2__sv2v_reg;
  assign r_9__1_ = r_9__1__sv2v_reg;
  assign r_9__0_ = r_9__0__sv2v_reg;
  assign r_10__15_ = r_10__15__sv2v_reg;
  assign r_10__14_ = r_10__14__sv2v_reg;
  assign r_10__13_ = r_10__13__sv2v_reg;
  assign r_10__12_ = r_10__12__sv2v_reg;
  assign r_10__11_ = r_10__11__sv2v_reg;
  assign r_10__10_ = r_10__10__sv2v_reg;
  assign r_10__9_ = r_10__9__sv2v_reg;
  assign r_10__8_ = r_10__8__sv2v_reg;
  assign r_10__7_ = r_10__7__sv2v_reg;
  assign r_10__6_ = r_10__6__sv2v_reg;
  assign r_10__5_ = r_10__5__sv2v_reg;
  assign r_10__4_ = r_10__4__sv2v_reg;
  assign r_10__3_ = r_10__3__sv2v_reg;
  assign r_10__2_ = r_10__2__sv2v_reg;
  assign r_10__1_ = r_10__1__sv2v_reg;
  assign r_10__0_ = r_10__0__sv2v_reg;
  assign r_11__15_ = r_11__15__sv2v_reg;
  assign r_11__14_ = r_11__14__sv2v_reg;
  assign r_11__13_ = r_11__13__sv2v_reg;
  assign r_11__12_ = r_11__12__sv2v_reg;
  assign r_11__11_ = r_11__11__sv2v_reg;
  assign r_11__10_ = r_11__10__sv2v_reg;
  assign r_11__9_ = r_11__9__sv2v_reg;
  assign r_11__8_ = r_11__8__sv2v_reg;
  assign r_11__7_ = r_11__7__sv2v_reg;
  assign r_11__6_ = r_11__6__sv2v_reg;
  assign r_11__5_ = r_11__5__sv2v_reg;
  assign r_11__4_ = r_11__4__sv2v_reg;
  assign r_11__3_ = r_11__3__sv2v_reg;
  assign r_11__2_ = r_11__2__sv2v_reg;
  assign r_11__1_ = r_11__1__sv2v_reg;
  assign r_11__0_ = r_11__0__sv2v_reg;
  assign r_12__15_ = r_12__15__sv2v_reg;
  assign r_12__14_ = r_12__14__sv2v_reg;
  assign r_12__13_ = r_12__13__sv2v_reg;
  assign r_12__12_ = r_12__12__sv2v_reg;
  assign r_12__11_ = r_12__11__sv2v_reg;
  assign r_12__10_ = r_12__10__sv2v_reg;
  assign r_12__9_ = r_12__9__sv2v_reg;
  assign r_12__8_ = r_12__8__sv2v_reg;
  assign r_12__7_ = r_12__7__sv2v_reg;
  assign r_12__6_ = r_12__6__sv2v_reg;
  assign r_12__5_ = r_12__5__sv2v_reg;
  assign r_12__4_ = r_12__4__sv2v_reg;
  assign r_12__3_ = r_12__3__sv2v_reg;
  assign r_12__2_ = r_12__2__sv2v_reg;
  assign r_12__1_ = r_12__1__sv2v_reg;
  assign r_12__0_ = r_12__0__sv2v_reg;
  assign r_13__15_ = r_13__15__sv2v_reg;
  assign r_13__14_ = r_13__14__sv2v_reg;
  assign r_13__13_ = r_13__13__sv2v_reg;
  assign r_13__12_ = r_13__12__sv2v_reg;
  assign r_13__11_ = r_13__11__sv2v_reg;
  assign r_13__10_ = r_13__10__sv2v_reg;
  assign r_13__9_ = r_13__9__sv2v_reg;
  assign r_13__8_ = r_13__8__sv2v_reg;
  assign r_13__7_ = r_13__7__sv2v_reg;
  assign r_13__6_ = r_13__6__sv2v_reg;
  assign r_13__5_ = r_13__5__sv2v_reg;
  assign r_13__4_ = r_13__4__sv2v_reg;
  assign r_13__3_ = r_13__3__sv2v_reg;
  assign r_13__2_ = r_13__2__sv2v_reg;
  assign r_13__1_ = r_13__1__sv2v_reg;
  assign r_13__0_ = r_13__0__sv2v_reg;
  assign r_14__15_ = r_14__15__sv2v_reg;
  assign r_14__14_ = r_14__14__sv2v_reg;
  assign r_14__13_ = r_14__13__sv2v_reg;
  assign r_14__12_ = r_14__12__sv2v_reg;
  assign r_14__11_ = r_14__11__sv2v_reg;
  assign r_14__10_ = r_14__10__sv2v_reg;
  assign r_14__9_ = r_14__9__sv2v_reg;
  assign r_14__8_ = r_14__8__sv2v_reg;
  assign r_14__7_ = r_14__7__sv2v_reg;
  assign r_14__6_ = r_14__6__sv2v_reg;
  assign r_14__5_ = r_14__5__sv2v_reg;
  assign r_14__4_ = r_14__4__sv2v_reg;
  assign r_14__3_ = r_14__3__sv2v_reg;
  assign r_14__2_ = r_14__2__sv2v_reg;
  assign r_14__1_ = r_14__1__sv2v_reg;
  assign r_14__0_ = r_14__0__sv2v_reg;
  assign r_15__15_ = r_15__15__sv2v_reg;
  assign r_15__14_ = r_15__14__sv2v_reg;
  assign r_15__13_ = r_15__13__sv2v_reg;
  assign r_15__12_ = r_15__12__sv2v_reg;
  assign r_15__11_ = r_15__11__sv2v_reg;
  assign r_15__10_ = r_15__10__sv2v_reg;
  assign r_15__9_ = r_15__9__sv2v_reg;
  assign r_15__8_ = r_15__8__sv2v_reg;
  assign r_15__7_ = r_15__7__sv2v_reg;
  assign r_15__6_ = r_15__6__sv2v_reg;
  assign r_15__5_ = r_15__5__sv2v_reg;
  assign r_15__4_ = r_15__4__sv2v_reg;
  assign r_15__3_ = r_15__3__sv2v_reg;
  assign r_15__2_ = r_15__2__sv2v_reg;
  assign r_15__1_ = r_15__1__sv2v_reg;
  assign r_15__0_ = r_15__0__sv2v_reg;
  assign r_16__15_ = r_16__15__sv2v_reg;
  assign r_16__14_ = r_16__14__sv2v_reg;
  assign r_16__13_ = r_16__13__sv2v_reg;
  assign r_16__12_ = r_16__12__sv2v_reg;
  assign r_16__11_ = r_16__11__sv2v_reg;
  assign r_16__10_ = r_16__10__sv2v_reg;
  assign r_16__9_ = r_16__9__sv2v_reg;
  assign r_16__8_ = r_16__8__sv2v_reg;
  assign r_16__7_ = r_16__7__sv2v_reg;
  assign r_16__6_ = r_16__6__sv2v_reg;
  assign r_16__5_ = r_16__5__sv2v_reg;
  assign r_16__4_ = r_16__4__sv2v_reg;
  assign r_16__3_ = r_16__3__sv2v_reg;
  assign r_16__2_ = r_16__2__sv2v_reg;
  assign r_16__1_ = r_16__1__sv2v_reg;
  assign r_16__0_ = r_16__0__sv2v_reg;
  assign r_17__15_ = r_17__15__sv2v_reg;
  assign r_17__14_ = r_17__14__sv2v_reg;
  assign r_17__13_ = r_17__13__sv2v_reg;
  assign r_17__12_ = r_17__12__sv2v_reg;
  assign r_17__11_ = r_17__11__sv2v_reg;
  assign r_17__10_ = r_17__10__sv2v_reg;
  assign r_17__9_ = r_17__9__sv2v_reg;
  assign r_17__8_ = r_17__8__sv2v_reg;
  assign r_17__7_ = r_17__7__sv2v_reg;
  assign r_17__6_ = r_17__6__sv2v_reg;
  assign r_17__5_ = r_17__5__sv2v_reg;
  assign r_17__4_ = r_17__4__sv2v_reg;
  assign r_17__3_ = r_17__3__sv2v_reg;
  assign r_17__2_ = r_17__2__sv2v_reg;
  assign r_17__1_ = r_17__1__sv2v_reg;
  assign r_17__0_ = r_17__0__sv2v_reg;
  assign r_18__15_ = r_18__15__sv2v_reg;
  assign r_18__14_ = r_18__14__sv2v_reg;
  assign r_18__13_ = r_18__13__sv2v_reg;
  assign r_18__12_ = r_18__12__sv2v_reg;
  assign r_18__11_ = r_18__11__sv2v_reg;
  assign r_18__10_ = r_18__10__sv2v_reg;
  assign r_18__9_ = r_18__9__sv2v_reg;
  assign r_18__8_ = r_18__8__sv2v_reg;
  assign r_18__7_ = r_18__7__sv2v_reg;
  assign r_18__6_ = r_18__6__sv2v_reg;
  assign r_18__5_ = r_18__5__sv2v_reg;
  assign r_18__4_ = r_18__4__sv2v_reg;
  assign r_18__3_ = r_18__3__sv2v_reg;
  assign r_18__2_ = r_18__2__sv2v_reg;
  assign r_18__1_ = r_18__1__sv2v_reg;
  assign r_18__0_ = r_18__0__sv2v_reg;
  assign r_19__15_ = r_19__15__sv2v_reg;
  assign r_19__14_ = r_19__14__sv2v_reg;
  assign r_19__13_ = r_19__13__sv2v_reg;
  assign r_19__12_ = r_19__12__sv2v_reg;
  assign r_19__11_ = r_19__11__sv2v_reg;
  assign r_19__10_ = r_19__10__sv2v_reg;
  assign r_19__9_ = r_19__9__sv2v_reg;
  assign r_19__8_ = r_19__8__sv2v_reg;
  assign r_19__7_ = r_19__7__sv2v_reg;
  assign r_19__6_ = r_19__6__sv2v_reg;
  assign r_19__5_ = r_19__5__sv2v_reg;
  assign r_19__4_ = r_19__4__sv2v_reg;
  assign r_19__3_ = r_19__3__sv2v_reg;
  assign r_19__2_ = r_19__2__sv2v_reg;
  assign r_19__1_ = r_19__1__sv2v_reg;
  assign r_19__0_ = r_19__0__sv2v_reg;
  assign r_20__15_ = r_20__15__sv2v_reg;
  assign r_20__14_ = r_20__14__sv2v_reg;
  assign r_20__13_ = r_20__13__sv2v_reg;
  assign r_20__12_ = r_20__12__sv2v_reg;
  assign r_20__11_ = r_20__11__sv2v_reg;
  assign r_20__10_ = r_20__10__sv2v_reg;
  assign r_20__9_ = r_20__9__sv2v_reg;
  assign r_20__8_ = r_20__8__sv2v_reg;
  assign r_20__7_ = r_20__7__sv2v_reg;
  assign r_20__6_ = r_20__6__sv2v_reg;
  assign r_20__5_ = r_20__5__sv2v_reg;
  assign r_20__4_ = r_20__4__sv2v_reg;
  assign r_20__3_ = r_20__3__sv2v_reg;
  assign r_20__2_ = r_20__2__sv2v_reg;
  assign r_20__1_ = r_20__1__sv2v_reg;
  assign r_20__0_ = r_20__0__sv2v_reg;
  assign r_21__15_ = r_21__15__sv2v_reg;
  assign r_21__14_ = r_21__14__sv2v_reg;
  assign r_21__13_ = r_21__13__sv2v_reg;
  assign r_21__12_ = r_21__12__sv2v_reg;
  assign r_21__11_ = r_21__11__sv2v_reg;
  assign r_21__10_ = r_21__10__sv2v_reg;
  assign r_21__9_ = r_21__9__sv2v_reg;
  assign r_21__8_ = r_21__8__sv2v_reg;
  assign r_21__7_ = r_21__7__sv2v_reg;
  assign r_21__6_ = r_21__6__sv2v_reg;
  assign r_21__5_ = r_21__5__sv2v_reg;
  assign r_21__4_ = r_21__4__sv2v_reg;
  assign r_21__3_ = r_21__3__sv2v_reg;
  assign r_21__2_ = r_21__2__sv2v_reg;
  assign r_21__1_ = r_21__1__sv2v_reg;
  assign r_21__0_ = r_21__0__sv2v_reg;
  assign r_22__15_ = r_22__15__sv2v_reg;
  assign r_22__14_ = r_22__14__sv2v_reg;
  assign r_22__13_ = r_22__13__sv2v_reg;
  assign r_22__12_ = r_22__12__sv2v_reg;
  assign r_22__11_ = r_22__11__sv2v_reg;
  assign r_22__10_ = r_22__10__sv2v_reg;
  assign r_22__9_ = r_22__9__sv2v_reg;
  assign r_22__8_ = r_22__8__sv2v_reg;
  assign r_22__7_ = r_22__7__sv2v_reg;
  assign r_22__6_ = r_22__6__sv2v_reg;
  assign r_22__5_ = r_22__5__sv2v_reg;
  assign r_22__4_ = r_22__4__sv2v_reg;
  assign r_22__3_ = r_22__3__sv2v_reg;
  assign r_22__2_ = r_22__2__sv2v_reg;
  assign r_22__1_ = r_22__1__sv2v_reg;
  assign r_22__0_ = r_22__0__sv2v_reg;
  assign r_23__15_ = r_23__15__sv2v_reg;
  assign r_23__14_ = r_23__14__sv2v_reg;
  assign r_23__13_ = r_23__13__sv2v_reg;
  assign r_23__12_ = r_23__12__sv2v_reg;
  assign r_23__11_ = r_23__11__sv2v_reg;
  assign r_23__10_ = r_23__10__sv2v_reg;
  assign r_23__9_ = r_23__9__sv2v_reg;
  assign r_23__8_ = r_23__8__sv2v_reg;
  assign r_23__7_ = r_23__7__sv2v_reg;
  assign r_23__6_ = r_23__6__sv2v_reg;
  assign r_23__5_ = r_23__5__sv2v_reg;
  assign r_23__4_ = r_23__4__sv2v_reg;
  assign r_23__3_ = r_23__3__sv2v_reg;
  assign r_23__2_ = r_23__2__sv2v_reg;
  assign r_23__1_ = r_23__1__sv2v_reg;
  assign r_23__0_ = r_23__0__sv2v_reg;
  assign r_24__15_ = r_24__15__sv2v_reg;
  assign r_24__14_ = r_24__14__sv2v_reg;
  assign r_24__13_ = r_24__13__sv2v_reg;
  assign r_24__12_ = r_24__12__sv2v_reg;
  assign r_24__11_ = r_24__11__sv2v_reg;
  assign r_24__10_ = r_24__10__sv2v_reg;
  assign r_24__9_ = r_24__9__sv2v_reg;
  assign r_24__8_ = r_24__8__sv2v_reg;
  assign r_24__7_ = r_24__7__sv2v_reg;
  assign r_24__6_ = r_24__6__sv2v_reg;
  assign r_24__5_ = r_24__5__sv2v_reg;
  assign r_24__4_ = r_24__4__sv2v_reg;
  assign r_24__3_ = r_24__3__sv2v_reg;
  assign r_24__2_ = r_24__2__sv2v_reg;
  assign r_24__1_ = r_24__1__sv2v_reg;
  assign r_24__0_ = r_24__0__sv2v_reg;
  assign r_25__15_ = r_25__15__sv2v_reg;
  assign r_25__14_ = r_25__14__sv2v_reg;
  assign r_25__13_ = r_25__13__sv2v_reg;
  assign r_25__12_ = r_25__12__sv2v_reg;
  assign r_25__11_ = r_25__11__sv2v_reg;
  assign r_25__10_ = r_25__10__sv2v_reg;
  assign r_25__9_ = r_25__9__sv2v_reg;
  assign r_25__8_ = r_25__8__sv2v_reg;
  assign r_25__7_ = r_25__7__sv2v_reg;
  assign r_25__6_ = r_25__6__sv2v_reg;
  assign r_25__5_ = r_25__5__sv2v_reg;
  assign r_25__4_ = r_25__4__sv2v_reg;
  assign r_25__3_ = r_25__3__sv2v_reg;
  assign r_25__2_ = r_25__2__sv2v_reg;
  assign r_25__1_ = r_25__1__sv2v_reg;
  assign r_25__0_ = r_25__0__sv2v_reg;
  assign r_26__15_ = r_26__15__sv2v_reg;
  assign r_26__14_ = r_26__14__sv2v_reg;
  assign r_26__13_ = r_26__13__sv2v_reg;
  assign r_26__12_ = r_26__12__sv2v_reg;
  assign r_26__11_ = r_26__11__sv2v_reg;
  assign r_26__10_ = r_26__10__sv2v_reg;
  assign r_26__9_ = r_26__9__sv2v_reg;
  assign r_26__8_ = r_26__8__sv2v_reg;
  assign r_26__7_ = r_26__7__sv2v_reg;
  assign r_26__6_ = r_26__6__sv2v_reg;
  assign r_26__5_ = r_26__5__sv2v_reg;
  assign r_26__4_ = r_26__4__sv2v_reg;
  assign r_26__3_ = r_26__3__sv2v_reg;
  assign r_26__2_ = r_26__2__sv2v_reg;
  assign r_26__1_ = r_26__1__sv2v_reg;
  assign r_26__0_ = r_26__0__sv2v_reg;
  assign r_27__15_ = r_27__15__sv2v_reg;
  assign r_27__14_ = r_27__14__sv2v_reg;
  assign r_27__13_ = r_27__13__sv2v_reg;
  assign r_27__12_ = r_27__12__sv2v_reg;
  assign r_27__11_ = r_27__11__sv2v_reg;
  assign r_27__10_ = r_27__10__sv2v_reg;
  assign r_27__9_ = r_27__9__sv2v_reg;
  assign r_27__8_ = r_27__8__sv2v_reg;
  assign r_27__7_ = r_27__7__sv2v_reg;
  assign r_27__6_ = r_27__6__sv2v_reg;
  assign r_27__5_ = r_27__5__sv2v_reg;
  assign r_27__4_ = r_27__4__sv2v_reg;
  assign r_27__3_ = r_27__3__sv2v_reg;
  assign r_27__2_ = r_27__2__sv2v_reg;
  assign r_27__1_ = r_27__1__sv2v_reg;
  assign r_27__0_ = r_27__0__sv2v_reg;
  assign r_28__15_ = r_28__15__sv2v_reg;
  assign r_28__14_ = r_28__14__sv2v_reg;
  assign r_28__13_ = r_28__13__sv2v_reg;
  assign r_28__12_ = r_28__12__sv2v_reg;
  assign r_28__11_ = r_28__11__sv2v_reg;
  assign r_28__10_ = r_28__10__sv2v_reg;
  assign r_28__9_ = r_28__9__sv2v_reg;
  assign r_28__8_ = r_28__8__sv2v_reg;
  assign r_28__7_ = r_28__7__sv2v_reg;
  assign r_28__6_ = r_28__6__sv2v_reg;
  assign r_28__5_ = r_28__5__sv2v_reg;
  assign r_28__4_ = r_28__4__sv2v_reg;
  assign r_28__3_ = r_28__3__sv2v_reg;
  assign r_28__2_ = r_28__2__sv2v_reg;
  assign r_28__1_ = r_28__1__sv2v_reg;
  assign r_28__0_ = r_28__0__sv2v_reg;
  assign r_29__15_ = r_29__15__sv2v_reg;
  assign r_29__14_ = r_29__14__sv2v_reg;
  assign r_29__13_ = r_29__13__sv2v_reg;
  assign r_29__12_ = r_29__12__sv2v_reg;
  assign r_29__11_ = r_29__11__sv2v_reg;
  assign r_29__10_ = r_29__10__sv2v_reg;
  assign r_29__9_ = r_29__9__sv2v_reg;
  assign r_29__8_ = r_29__8__sv2v_reg;
  assign r_29__7_ = r_29__7__sv2v_reg;
  assign r_29__6_ = r_29__6__sv2v_reg;
  assign r_29__5_ = r_29__5__sv2v_reg;
  assign r_29__4_ = r_29__4__sv2v_reg;
  assign r_29__3_ = r_29__3__sv2v_reg;
  assign r_29__2_ = r_29__2__sv2v_reg;
  assign r_29__1_ = r_29__1__sv2v_reg;
  assign r_29__0_ = r_29__0__sv2v_reg;
  assign r_30__15_ = r_30__15__sv2v_reg;
  assign r_30__14_ = r_30__14__sv2v_reg;
  assign r_30__13_ = r_30__13__sv2v_reg;
  assign r_30__12_ = r_30__12__sv2v_reg;
  assign r_30__11_ = r_30__11__sv2v_reg;
  assign r_30__10_ = r_30__10__sv2v_reg;
  assign r_30__9_ = r_30__9__sv2v_reg;
  assign r_30__8_ = r_30__8__sv2v_reg;
  assign r_30__7_ = r_30__7__sv2v_reg;
  assign r_30__6_ = r_30__6__sv2v_reg;
  assign r_30__5_ = r_30__5__sv2v_reg;
  assign r_30__4_ = r_30__4__sv2v_reg;
  assign r_30__3_ = r_30__3__sv2v_reg;
  assign r_30__2_ = r_30__2__sv2v_reg;
  assign r_30__1_ = r_30__1__sv2v_reg;
  assign r_30__0_ = r_30__0__sv2v_reg;
  assign r_31__15_ = r_31__15__sv2v_reg;
  assign r_31__14_ = r_31__14__sv2v_reg;
  assign r_31__13_ = r_31__13__sv2v_reg;
  assign r_31__12_ = r_31__12__sv2v_reg;
  assign r_31__11_ = r_31__11__sv2v_reg;
  assign r_31__10_ = r_31__10__sv2v_reg;
  assign r_31__9_ = r_31__9__sv2v_reg;
  assign r_31__8_ = r_31__8__sv2v_reg;
  assign r_31__7_ = r_31__7__sv2v_reg;
  assign r_31__6_ = r_31__6__sv2v_reg;
  assign r_31__5_ = r_31__5__sv2v_reg;
  assign r_31__4_ = r_31__4__sv2v_reg;
  assign r_31__3_ = r_31__3__sv2v_reg;
  assign r_31__2_ = r_31__2__sv2v_reg;
  assign r_31__1_ = r_31__1__sv2v_reg;
  assign r_31__0_ = r_31__0__sv2v_reg;
  assign N62 = sel_i[1] & sel_i[0];
  assign N64 = N63 & N66;
  assign N67 = sel_i[3] & sel_i[2];
  assign N69 = N68 & N71;
  assign N72 = sel_i[5] & sel_i[4];
  assign N74 = N73 & N76;
  assign N77 = sel_i[7] & sel_i[6];
  assign N79 = N78 & N81;
  assign N82 = sel_i[9] & sel_i[8];
  assign N84 = N83 & N86;
  assign N87 = sel_i[11] & sel_i[10];
  assign N89 = N88 & N91;
  assign N92 = sel_i[13] & sel_i[12];
  assign N94 = N93 & N96;
  assign N97 = sel_i[15] & sel_i[14];
  assign N99 = N98 & N101;
  assign N102 = sel_i[17] & sel_i[16];
  assign N104 = N103 & N106;
  assign N107 = sel_i[19] & sel_i[18];
  assign N109 = N108 & N111;
  assign N112 = sel_i[21] & sel_i[20];
  assign N114 = N113 & N116;
  assign N117 = sel_i[23] & sel_i[22];
  assign N119 = N118 & N121;
  assign N122 = sel_i[25] & sel_i[24];
  assign N124 = N123 & N126;
  assign N127 = sel_i[27] & sel_i[26];
  assign N129 = N128 & N131;
  assign N132 = sel_i[29] & sel_i[28];
  assign N134 = N133 & N136;
  assign N137 = sel_i[31] & sel_i[30];
  assign N139 = N138 & N141;
  assign N142 = sel_i[33] & sel_i[32];
  assign N144 = N143 & N146;
  assign N147 = sel_i[35] & sel_i[34];
  assign N149 = N148 & N151;
  assign N152 = sel_i[37] & sel_i[36];
  assign N154 = N153 & N156;
  assign N157 = sel_i[39] & sel_i[38];
  assign N159 = N158 & N161;
  assign N162 = sel_i[41] & sel_i[40];
  assign N164 = N163 & N166;
  assign N167 = sel_i[43] & sel_i[42];
  assign N169 = N168 & N171;
  assign N172 = sel_i[45] & sel_i[44];
  assign N174 = N173 & N176;
  assign N177 = sel_i[47] & sel_i[46];
  assign N179 = N178 & N181;
  assign N182 = sel_i[49] & sel_i[48];
  assign N184 = N183 & N186;
  assign N187 = sel_i[51] & sel_i[50];
  assign N189 = N188 & N191;
  assign N192 = sel_i[53] & sel_i[52];
  assign N194 = N193 & N196;
  assign N197 = sel_i[55] & sel_i[54];
  assign N199 = N198 & N201;
  assign N202 = sel_i[57] & sel_i[56];
  assign N204 = N203 & N206;
  assign N207 = sel_i[59] & sel_i[58];
  assign N209 = N208 & N211;
  assign N212 = sel_i[61] & sel_i[60];
  assign N214 = N213 & N216;
  assign N218 = sel_i[63] | N217;
  assign N220 = sel_i[63] & sel_i[62];
  assign N222 = N221 & N217;
  assign N66 = ~sel_i[0];
  assign N71 = ~sel_i[2];
  assign N76 = ~sel_i[4];
  assign N81 = ~sel_i[6];
  assign N86 = ~sel_i[8];
  assign N91 = ~sel_i[10];
  assign N96 = ~sel_i[12];
  assign N101 = ~sel_i[14];
  assign N106 = ~sel_i[16];
  assign N111 = ~sel_i[18];
  assign N116 = ~sel_i[20];
  assign N121 = ~sel_i[22];
  assign N126 = ~sel_i[24];
  assign N131 = ~sel_i[26];
  assign N136 = ~sel_i[28];
  assign N141 = ~sel_i[30];
  assign N146 = ~sel_i[32];
  assign N151 = ~sel_i[34];
  assign N156 = ~sel_i[36];
  assign N161 = ~sel_i[38];
  assign N166 = ~sel_i[40];
  assign N171 = ~sel_i[42];
  assign N176 = ~sel_i[44];
  assign N181 = ~sel_i[46];
  assign N186 = ~sel_i[48];
  assign N191 = ~sel_i[50];
  assign N196 = ~sel_i[52];
  assign N201 = ~sel_i[54];
  assign N206 = ~sel_i[56];
  assign N211 = ~sel_i[58];
  assign N216 = ~sel_i[60];
  assign { r_n_0__15_, r_n_0__14_, r_n_0__13_, r_n_0__12_, r_n_0__11_, r_n_0__10_, r_n_0__9_, r_n_0__8_, r_n_0__7_, r_n_0__6_, r_n_0__5_, r_n_0__4_, r_n_0__3_, r_n_0__2_, r_n_0__1_, r_n_0__0_ } = (N0)? { r_1__15_, r_1__14_, r_1__13_, r_1__12_, r_1__11_, r_1__10_, r_1__9_, r_1__8_, r_1__7_, r_1__6_, r_1__5_, r_1__4_, r_1__3_, r_1__2_, r_1__1_, r_1__0_ } : 
                                                                                                                                                                                                    (N1)? data_i : 1'b0;
  assign N0 = sel_i[0];
  assign N1 = N66;
  assign { r_n_1__15_, r_n_1__14_, r_n_1__13_, r_n_1__12_, r_n_1__11_, r_n_1__10_, r_n_1__9_, r_n_1__8_, r_n_1__7_, r_n_1__6_, r_n_1__5_, r_n_1__4_, r_n_1__3_, r_n_1__2_, r_n_1__1_, r_n_1__0_ } = (N2)? { r_2__15_, r_2__14_, r_2__13_, r_2__12_, r_2__11_, r_2__10_, r_2__9_, r_2__8_, r_2__7_, r_2__6_, r_2__5_, r_2__4_, r_2__3_, r_2__2_, r_2__1_, r_2__0_ } : 
                                                                                                                                                                                                    (N3)? data_i : 1'b0;
  assign N2 = sel_i[2];
  assign N3 = N71;
  assign { r_n_2__15_, r_n_2__14_, r_n_2__13_, r_n_2__12_, r_n_2__11_, r_n_2__10_, r_n_2__9_, r_n_2__8_, r_n_2__7_, r_n_2__6_, r_n_2__5_, r_n_2__4_, r_n_2__3_, r_n_2__2_, r_n_2__1_, r_n_2__0_ } = (N4)? { r_3__15_, r_3__14_, r_3__13_, r_3__12_, r_3__11_, r_3__10_, r_3__9_, r_3__8_, r_3__7_, r_3__6_, r_3__5_, r_3__4_, r_3__3_, r_3__2_, r_3__1_, r_3__0_ } : 
                                                                                                                                                                                                    (N5)? data_i : 1'b0;
  assign N4 = sel_i[4];
  assign N5 = N76;
  assign { r_n_3__15_, r_n_3__14_, r_n_3__13_, r_n_3__12_, r_n_3__11_, r_n_3__10_, r_n_3__9_, r_n_3__8_, r_n_3__7_, r_n_3__6_, r_n_3__5_, r_n_3__4_, r_n_3__3_, r_n_3__2_, r_n_3__1_, r_n_3__0_ } = (N6)? { r_4__15_, r_4__14_, r_4__13_, r_4__12_, r_4__11_, r_4__10_, r_4__9_, r_4__8_, r_4__7_, r_4__6_, r_4__5_, r_4__4_, r_4__3_, r_4__2_, r_4__1_, r_4__0_ } : 
                                                                                                                                                                                                    (N7)? data_i : 1'b0;
  assign N6 = sel_i[6];
  assign N7 = N81;
  assign { r_n_4__15_, r_n_4__14_, r_n_4__13_, r_n_4__12_, r_n_4__11_, r_n_4__10_, r_n_4__9_, r_n_4__8_, r_n_4__7_, r_n_4__6_, r_n_4__5_, r_n_4__4_, r_n_4__3_, r_n_4__2_, r_n_4__1_, r_n_4__0_ } = (N8)? { r_5__15_, r_5__14_, r_5__13_, r_5__12_, r_5__11_, r_5__10_, r_5__9_, r_5__8_, r_5__7_, r_5__6_, r_5__5_, r_5__4_, r_5__3_, r_5__2_, r_5__1_, r_5__0_ } : 
                                                                                                                                                                                                    (N9)? data_i : 1'b0;
  assign N8 = sel_i[8];
  assign N9 = N86;
  assign { r_n_5__15_, r_n_5__14_, r_n_5__13_, r_n_5__12_, r_n_5__11_, r_n_5__10_, r_n_5__9_, r_n_5__8_, r_n_5__7_, r_n_5__6_, r_n_5__5_, r_n_5__4_, r_n_5__3_, r_n_5__2_, r_n_5__1_, r_n_5__0_ } = (N10)? { r_6__15_, r_6__14_, r_6__13_, r_6__12_, r_6__11_, r_6__10_, r_6__9_, r_6__8_, r_6__7_, r_6__6_, r_6__5_, r_6__4_, r_6__3_, r_6__2_, r_6__1_, r_6__0_ } : 
                                                                                                                                                                                                    (N11)? data_i : 1'b0;
  assign N10 = sel_i[10];
  assign N11 = N91;
  assign { r_n_6__15_, r_n_6__14_, r_n_6__13_, r_n_6__12_, r_n_6__11_, r_n_6__10_, r_n_6__9_, r_n_6__8_, r_n_6__7_, r_n_6__6_, r_n_6__5_, r_n_6__4_, r_n_6__3_, r_n_6__2_, r_n_6__1_, r_n_6__0_ } = (N12)? { r_7__15_, r_7__14_, r_7__13_, r_7__12_, r_7__11_, r_7__10_, r_7__9_, r_7__8_, r_7__7_, r_7__6_, r_7__5_, r_7__4_, r_7__3_, r_7__2_, r_7__1_, r_7__0_ } : 
                                                                                                                                                                                                    (N13)? data_i : 1'b0;
  assign N12 = sel_i[12];
  assign N13 = N96;
  assign { r_n_7__15_, r_n_7__14_, r_n_7__13_, r_n_7__12_, r_n_7__11_, r_n_7__10_, r_n_7__9_, r_n_7__8_, r_n_7__7_, r_n_7__6_, r_n_7__5_, r_n_7__4_, r_n_7__3_, r_n_7__2_, r_n_7__1_, r_n_7__0_ } = (N14)? { r_8__15_, r_8__14_, r_8__13_, r_8__12_, r_8__11_, r_8__10_, r_8__9_, r_8__8_, r_8__7_, r_8__6_, r_8__5_, r_8__4_, r_8__3_, r_8__2_, r_8__1_, r_8__0_ } : 
                                                                                                                                                                                                    (N15)? data_i : 1'b0;
  assign N14 = sel_i[14];
  assign N15 = N101;
  assign { r_n_8__15_, r_n_8__14_, r_n_8__13_, r_n_8__12_, r_n_8__11_, r_n_8__10_, r_n_8__9_, r_n_8__8_, r_n_8__7_, r_n_8__6_, r_n_8__5_, r_n_8__4_, r_n_8__3_, r_n_8__2_, r_n_8__1_, r_n_8__0_ } = (N16)? { r_9__15_, r_9__14_, r_9__13_, r_9__12_, r_9__11_, r_9__10_, r_9__9_, r_9__8_, r_9__7_, r_9__6_, r_9__5_, r_9__4_, r_9__3_, r_9__2_, r_9__1_, r_9__0_ } : 
                                                                                                                                                                                                    (N17)? data_i : 1'b0;
  assign N16 = sel_i[16];
  assign N17 = N106;
  assign { r_n_9__15_, r_n_9__14_, r_n_9__13_, r_n_9__12_, r_n_9__11_, r_n_9__10_, r_n_9__9_, r_n_9__8_, r_n_9__7_, r_n_9__6_, r_n_9__5_, r_n_9__4_, r_n_9__3_, r_n_9__2_, r_n_9__1_, r_n_9__0_ } = (N18)? { r_10__15_, r_10__14_, r_10__13_, r_10__12_, r_10__11_, r_10__10_, r_10__9_, r_10__8_, r_10__7_, r_10__6_, r_10__5_, r_10__4_, r_10__3_, r_10__2_, r_10__1_, r_10__0_ } : 
                                                                                                                                                                                                    (N19)? data_i : 1'b0;
  assign N18 = sel_i[18];
  assign N19 = N111;
  assign { r_n_10__15_, r_n_10__14_, r_n_10__13_, r_n_10__12_, r_n_10__11_, r_n_10__10_, r_n_10__9_, r_n_10__8_, r_n_10__7_, r_n_10__6_, r_n_10__5_, r_n_10__4_, r_n_10__3_, r_n_10__2_, r_n_10__1_, r_n_10__0_ } = (N20)? { r_11__15_, r_11__14_, r_11__13_, r_11__12_, r_11__11_, r_11__10_, r_11__9_, r_11__8_, r_11__7_, r_11__6_, r_11__5_, r_11__4_, r_11__3_, r_11__2_, r_11__1_, r_11__0_ } : 
                                                                                                                                                                                                                    (N21)? data_i : 1'b0;
  assign N20 = sel_i[20];
  assign N21 = N116;
  assign { r_n_11__15_, r_n_11__14_, r_n_11__13_, r_n_11__12_, r_n_11__11_, r_n_11__10_, r_n_11__9_, r_n_11__8_, r_n_11__7_, r_n_11__6_, r_n_11__5_, r_n_11__4_, r_n_11__3_, r_n_11__2_, r_n_11__1_, r_n_11__0_ } = (N22)? { r_12__15_, r_12__14_, r_12__13_, r_12__12_, r_12__11_, r_12__10_, r_12__9_, r_12__8_, r_12__7_, r_12__6_, r_12__5_, r_12__4_, r_12__3_, r_12__2_, r_12__1_, r_12__0_ } : 
                                                                                                                                                                                                                    (N23)? data_i : 1'b0;
  assign N22 = sel_i[22];
  assign N23 = N121;
  assign { r_n_12__15_, r_n_12__14_, r_n_12__13_, r_n_12__12_, r_n_12__11_, r_n_12__10_, r_n_12__9_, r_n_12__8_, r_n_12__7_, r_n_12__6_, r_n_12__5_, r_n_12__4_, r_n_12__3_, r_n_12__2_, r_n_12__1_, r_n_12__0_ } = (N24)? { r_13__15_, r_13__14_, r_13__13_, r_13__12_, r_13__11_, r_13__10_, r_13__9_, r_13__8_, r_13__7_, r_13__6_, r_13__5_, r_13__4_, r_13__3_, r_13__2_, r_13__1_, r_13__0_ } : 
                                                                                                                                                                                                                    (N25)? data_i : 1'b0;
  assign N24 = sel_i[24];
  assign N25 = N126;
  assign { r_n_13__15_, r_n_13__14_, r_n_13__13_, r_n_13__12_, r_n_13__11_, r_n_13__10_, r_n_13__9_, r_n_13__8_, r_n_13__7_, r_n_13__6_, r_n_13__5_, r_n_13__4_, r_n_13__3_, r_n_13__2_, r_n_13__1_, r_n_13__0_ } = (N26)? { r_14__15_, r_14__14_, r_14__13_, r_14__12_, r_14__11_, r_14__10_, r_14__9_, r_14__8_, r_14__7_, r_14__6_, r_14__5_, r_14__4_, r_14__3_, r_14__2_, r_14__1_, r_14__0_ } : 
                                                                                                                                                                                                                    (N27)? data_i : 1'b0;
  assign N26 = sel_i[26];
  assign N27 = N131;
  assign { r_n_14__15_, r_n_14__14_, r_n_14__13_, r_n_14__12_, r_n_14__11_, r_n_14__10_, r_n_14__9_, r_n_14__8_, r_n_14__7_, r_n_14__6_, r_n_14__5_, r_n_14__4_, r_n_14__3_, r_n_14__2_, r_n_14__1_, r_n_14__0_ } = (N28)? { r_15__15_, r_15__14_, r_15__13_, r_15__12_, r_15__11_, r_15__10_, r_15__9_, r_15__8_, r_15__7_, r_15__6_, r_15__5_, r_15__4_, r_15__3_, r_15__2_, r_15__1_, r_15__0_ } : 
                                                                                                                                                                                                                    (N29)? data_i : 1'b0;
  assign N28 = sel_i[28];
  assign N29 = N136;
  assign { r_n_15__15_, r_n_15__14_, r_n_15__13_, r_n_15__12_, r_n_15__11_, r_n_15__10_, r_n_15__9_, r_n_15__8_, r_n_15__7_, r_n_15__6_, r_n_15__5_, r_n_15__4_, r_n_15__3_, r_n_15__2_, r_n_15__1_, r_n_15__0_ } = (N30)? { r_16__15_, r_16__14_, r_16__13_, r_16__12_, r_16__11_, r_16__10_, r_16__9_, r_16__8_, r_16__7_, r_16__6_, r_16__5_, r_16__4_, r_16__3_, r_16__2_, r_16__1_, r_16__0_ } : 
                                                                                                                                                                                                                    (N31)? data_i : 1'b0;
  assign N30 = sel_i[30];
  assign N31 = N141;
  assign { r_n_16__15_, r_n_16__14_, r_n_16__13_, r_n_16__12_, r_n_16__11_, r_n_16__10_, r_n_16__9_, r_n_16__8_, r_n_16__7_, r_n_16__6_, r_n_16__5_, r_n_16__4_, r_n_16__3_, r_n_16__2_, r_n_16__1_, r_n_16__0_ } = (N32)? { r_17__15_, r_17__14_, r_17__13_, r_17__12_, r_17__11_, r_17__10_, r_17__9_, r_17__8_, r_17__7_, r_17__6_, r_17__5_, r_17__4_, r_17__3_, r_17__2_, r_17__1_, r_17__0_ } : 
                                                                                                                                                                                                                    (N33)? data_i : 1'b0;
  assign N32 = sel_i[32];
  assign N33 = N146;
  assign { r_n_17__15_, r_n_17__14_, r_n_17__13_, r_n_17__12_, r_n_17__11_, r_n_17__10_, r_n_17__9_, r_n_17__8_, r_n_17__7_, r_n_17__6_, r_n_17__5_, r_n_17__4_, r_n_17__3_, r_n_17__2_, r_n_17__1_, r_n_17__0_ } = (N34)? { r_18__15_, r_18__14_, r_18__13_, r_18__12_, r_18__11_, r_18__10_, r_18__9_, r_18__8_, r_18__7_, r_18__6_, r_18__5_, r_18__4_, r_18__3_, r_18__2_, r_18__1_, r_18__0_ } : 
                                                                                                                                                                                                                    (N35)? data_i : 1'b0;
  assign N34 = sel_i[34];
  assign N35 = N151;
  assign { r_n_18__15_, r_n_18__14_, r_n_18__13_, r_n_18__12_, r_n_18__11_, r_n_18__10_, r_n_18__9_, r_n_18__8_, r_n_18__7_, r_n_18__6_, r_n_18__5_, r_n_18__4_, r_n_18__3_, r_n_18__2_, r_n_18__1_, r_n_18__0_ } = (N36)? { r_19__15_, r_19__14_, r_19__13_, r_19__12_, r_19__11_, r_19__10_, r_19__9_, r_19__8_, r_19__7_, r_19__6_, r_19__5_, r_19__4_, r_19__3_, r_19__2_, r_19__1_, r_19__0_ } : 
                                                                                                                                                                                                                    (N37)? data_i : 1'b0;
  assign N36 = sel_i[36];
  assign N37 = N156;
  assign { r_n_19__15_, r_n_19__14_, r_n_19__13_, r_n_19__12_, r_n_19__11_, r_n_19__10_, r_n_19__9_, r_n_19__8_, r_n_19__7_, r_n_19__6_, r_n_19__5_, r_n_19__4_, r_n_19__3_, r_n_19__2_, r_n_19__1_, r_n_19__0_ } = (N38)? { r_20__15_, r_20__14_, r_20__13_, r_20__12_, r_20__11_, r_20__10_, r_20__9_, r_20__8_, r_20__7_, r_20__6_, r_20__5_, r_20__4_, r_20__3_, r_20__2_, r_20__1_, r_20__0_ } : 
                                                                                                                                                                                                                    (N39)? data_i : 1'b0;
  assign N38 = sel_i[38];
  assign N39 = N161;
  assign { r_n_20__15_, r_n_20__14_, r_n_20__13_, r_n_20__12_, r_n_20__11_, r_n_20__10_, r_n_20__9_, r_n_20__8_, r_n_20__7_, r_n_20__6_, r_n_20__5_, r_n_20__4_, r_n_20__3_, r_n_20__2_, r_n_20__1_, r_n_20__0_ } = (N40)? { r_21__15_, r_21__14_, r_21__13_, r_21__12_, r_21__11_, r_21__10_, r_21__9_, r_21__8_, r_21__7_, r_21__6_, r_21__5_, r_21__4_, r_21__3_, r_21__2_, r_21__1_, r_21__0_ } : 
                                                                                                                                                                                                                    (N41)? data_i : 1'b0;
  assign N40 = sel_i[40];
  assign N41 = N166;
  assign { r_n_21__15_, r_n_21__14_, r_n_21__13_, r_n_21__12_, r_n_21__11_, r_n_21__10_, r_n_21__9_, r_n_21__8_, r_n_21__7_, r_n_21__6_, r_n_21__5_, r_n_21__4_, r_n_21__3_, r_n_21__2_, r_n_21__1_, r_n_21__0_ } = (N42)? { r_22__15_, r_22__14_, r_22__13_, r_22__12_, r_22__11_, r_22__10_, r_22__9_, r_22__8_, r_22__7_, r_22__6_, r_22__5_, r_22__4_, r_22__3_, r_22__2_, r_22__1_, r_22__0_ } : 
                                                                                                                                                                                                                    (N43)? data_i : 1'b0;
  assign N42 = sel_i[42];
  assign N43 = N171;
  assign { r_n_22__15_, r_n_22__14_, r_n_22__13_, r_n_22__12_, r_n_22__11_, r_n_22__10_, r_n_22__9_, r_n_22__8_, r_n_22__7_, r_n_22__6_, r_n_22__5_, r_n_22__4_, r_n_22__3_, r_n_22__2_, r_n_22__1_, r_n_22__0_ } = (N44)? { r_23__15_, r_23__14_, r_23__13_, r_23__12_, r_23__11_, r_23__10_, r_23__9_, r_23__8_, r_23__7_, r_23__6_, r_23__5_, r_23__4_, r_23__3_, r_23__2_, r_23__1_, r_23__0_ } : 
                                                                                                                                                                                                                    (N45)? data_i : 1'b0;
  assign N44 = sel_i[44];
  assign N45 = N176;
  assign { r_n_23__15_, r_n_23__14_, r_n_23__13_, r_n_23__12_, r_n_23__11_, r_n_23__10_, r_n_23__9_, r_n_23__8_, r_n_23__7_, r_n_23__6_, r_n_23__5_, r_n_23__4_, r_n_23__3_, r_n_23__2_, r_n_23__1_, r_n_23__0_ } = (N46)? { r_24__15_, r_24__14_, r_24__13_, r_24__12_, r_24__11_, r_24__10_, r_24__9_, r_24__8_, r_24__7_, r_24__6_, r_24__5_, r_24__4_, r_24__3_, r_24__2_, r_24__1_, r_24__0_ } : 
                                                                                                                                                                                                                    (N47)? data_i : 1'b0;
  assign N46 = sel_i[46];
  assign N47 = N181;
  assign { r_n_24__15_, r_n_24__14_, r_n_24__13_, r_n_24__12_, r_n_24__11_, r_n_24__10_, r_n_24__9_, r_n_24__8_, r_n_24__7_, r_n_24__6_, r_n_24__5_, r_n_24__4_, r_n_24__3_, r_n_24__2_, r_n_24__1_, r_n_24__0_ } = (N48)? { r_25__15_, r_25__14_, r_25__13_, r_25__12_, r_25__11_, r_25__10_, r_25__9_, r_25__8_, r_25__7_, r_25__6_, r_25__5_, r_25__4_, r_25__3_, r_25__2_, r_25__1_, r_25__0_ } : 
                                                                                                                                                                                                                    (N49)? data_i : 1'b0;
  assign N48 = sel_i[48];
  assign N49 = N186;
  assign { r_n_25__15_, r_n_25__14_, r_n_25__13_, r_n_25__12_, r_n_25__11_, r_n_25__10_, r_n_25__9_, r_n_25__8_, r_n_25__7_, r_n_25__6_, r_n_25__5_, r_n_25__4_, r_n_25__3_, r_n_25__2_, r_n_25__1_, r_n_25__0_ } = (N50)? { r_26__15_, r_26__14_, r_26__13_, r_26__12_, r_26__11_, r_26__10_, r_26__9_, r_26__8_, r_26__7_, r_26__6_, r_26__5_, r_26__4_, r_26__3_, r_26__2_, r_26__1_, r_26__0_ } : 
                                                                                                                                                                                                                    (N51)? data_i : 1'b0;
  assign N50 = sel_i[50];
  assign N51 = N191;
  assign { r_n_26__15_, r_n_26__14_, r_n_26__13_, r_n_26__12_, r_n_26__11_, r_n_26__10_, r_n_26__9_, r_n_26__8_, r_n_26__7_, r_n_26__6_, r_n_26__5_, r_n_26__4_, r_n_26__3_, r_n_26__2_, r_n_26__1_, r_n_26__0_ } = (N52)? { r_27__15_, r_27__14_, r_27__13_, r_27__12_, r_27__11_, r_27__10_, r_27__9_, r_27__8_, r_27__7_, r_27__6_, r_27__5_, r_27__4_, r_27__3_, r_27__2_, r_27__1_, r_27__0_ } : 
                                                                                                                                                                                                                    (N53)? data_i : 1'b0;
  assign N52 = sel_i[52];
  assign N53 = N196;
  assign { r_n_27__15_, r_n_27__14_, r_n_27__13_, r_n_27__12_, r_n_27__11_, r_n_27__10_, r_n_27__9_, r_n_27__8_, r_n_27__7_, r_n_27__6_, r_n_27__5_, r_n_27__4_, r_n_27__3_, r_n_27__2_, r_n_27__1_, r_n_27__0_ } = (N54)? { r_28__15_, r_28__14_, r_28__13_, r_28__12_, r_28__11_, r_28__10_, r_28__9_, r_28__8_, r_28__7_, r_28__6_, r_28__5_, r_28__4_, r_28__3_, r_28__2_, r_28__1_, r_28__0_ } : 
                                                                                                                                                                                                                    (N55)? data_i : 1'b0;
  assign N54 = sel_i[54];
  assign N55 = N201;
  assign { r_n_28__15_, r_n_28__14_, r_n_28__13_, r_n_28__12_, r_n_28__11_, r_n_28__10_, r_n_28__9_, r_n_28__8_, r_n_28__7_, r_n_28__6_, r_n_28__5_, r_n_28__4_, r_n_28__3_, r_n_28__2_, r_n_28__1_, r_n_28__0_ } = (N56)? { r_29__15_, r_29__14_, r_29__13_, r_29__12_, r_29__11_, r_29__10_, r_29__9_, r_29__8_, r_29__7_, r_29__6_, r_29__5_, r_29__4_, r_29__3_, r_29__2_, r_29__1_, r_29__0_ } : 
                                                                                                                                                                                                                    (N57)? data_i : 1'b0;
  assign N56 = sel_i[56];
  assign N57 = N206;
  assign { r_n_29__15_, r_n_29__14_, r_n_29__13_, r_n_29__12_, r_n_29__11_, r_n_29__10_, r_n_29__9_, r_n_29__8_, r_n_29__7_, r_n_29__6_, r_n_29__5_, r_n_29__4_, r_n_29__3_, r_n_29__2_, r_n_29__1_, r_n_29__0_ } = (N58)? { r_30__15_, r_30__14_, r_30__13_, r_30__12_, r_30__11_, r_30__10_, r_30__9_, r_30__8_, r_30__7_, r_30__6_, r_30__5_, r_30__4_, r_30__3_, r_30__2_, r_30__1_, r_30__0_ } : 
                                                                                                                                                                                                                    (N59)? data_i : 1'b0;
  assign N58 = sel_i[58];
  assign N59 = N211;
  assign { r_n_30__15_, r_n_30__14_, r_n_30__13_, r_n_30__12_, r_n_30__11_, r_n_30__10_, r_n_30__9_, r_n_30__8_, r_n_30__7_, r_n_30__6_, r_n_30__5_, r_n_30__4_, r_n_30__3_, r_n_30__2_, r_n_30__1_, r_n_30__0_ } = (N60)? { r_31__15_, r_31__14_, r_31__13_, r_31__12_, r_31__11_, r_31__10_, r_31__9_, r_31__8_, r_31__7_, r_31__6_, r_31__5_, r_31__4_, r_31__3_, r_31__2_, r_31__1_, r_31__0_ } : 
                                                                                                                                                                                                                    (N61)? data_i : 1'b0;
  assign N60 = sel_i[60];
  assign N61 = N216;
  assign N63 = ~sel_i[1];
  assign N65 = N62 | N64;
  assign N68 = ~sel_i[3];
  assign N70 = N67 | N69;
  assign N73 = ~sel_i[5];
  assign N75 = N72 | N74;
  assign N78 = ~sel_i[7];
  assign N80 = N77 | N79;
  assign N83 = ~sel_i[9];
  assign N85 = N82 | N84;
  assign N88 = ~sel_i[11];
  assign N90 = N87 | N89;
  assign N93 = ~sel_i[13];
  assign N95 = N92 | N94;
  assign N98 = ~sel_i[15];
  assign N100 = N97 | N99;
  assign N103 = ~sel_i[17];
  assign N105 = N102 | N104;
  assign N108 = ~sel_i[19];
  assign N110 = N107 | N109;
  assign N113 = ~sel_i[21];
  assign N115 = N112 | N114;
  assign N118 = ~sel_i[23];
  assign N120 = N117 | N119;
  assign N123 = ~sel_i[25];
  assign N125 = N122 | N124;
  assign N128 = ~sel_i[27];
  assign N130 = N127 | N129;
  assign N133 = ~sel_i[29];
  assign N135 = N132 | N134;
  assign N138 = ~sel_i[31];
  assign N140 = N137 | N139;
  assign N143 = ~sel_i[33];
  assign N145 = N142 | N144;
  assign N148 = ~sel_i[35];
  assign N150 = N147 | N149;
  assign N153 = ~sel_i[37];
  assign N155 = N152 | N154;
  assign N158 = ~sel_i[39];
  assign N160 = N157 | N159;
  assign N163 = ~sel_i[41];
  assign N165 = N162 | N164;
  assign N168 = ~sel_i[43];
  assign N170 = N167 | N169;
  assign N173 = ~sel_i[45];
  assign N175 = N172 | N174;
  assign N178 = ~sel_i[47];
  assign N180 = N177 | N179;
  assign N183 = ~sel_i[49];
  assign N185 = N182 | N184;
  assign N188 = ~sel_i[51];
  assign N190 = N187 | N189;
  assign N193 = ~sel_i[53];
  assign N195 = N192 | N194;
  assign N198 = ~sel_i[55];
  assign N200 = N197 | N199;
  assign N203 = ~sel_i[57];
  assign N205 = N202 | N204;
  assign N208 = ~sel_i[59];
  assign N210 = N207 | N209;
  assign N213 = ~sel_i[61];
  assign N215 = N212 | N214;
  assign N217 = ~sel_i[62];
  assign N219 = ~N218;
  assign N221 = ~sel_i[63];
  assign N223 = N220 | N222;
  assign N224 = ~N65;
  assign N225 = ~N70;
  assign N226 = ~N75;
  assign N227 = ~N80;
  assign N228 = ~N85;
  assign N229 = ~N90;
  assign N230 = ~N95;
  assign N231 = ~N100;
  assign N232 = ~N105;
  assign N233 = ~N110;
  assign N234 = ~N115;
  assign N235 = ~N120;
  assign N236 = ~N125;
  assign N237 = ~N130;
  assign N238 = ~N135;
  assign N239 = ~N140;
  assign N240 = ~N145;
  assign N241 = ~N150;
  assign N242 = ~N155;
  assign N243 = ~N160;
  assign N244 = ~N165;
  assign N245 = ~N170;
  assign N246 = ~N175;
  assign N247 = ~N180;
  assign N248 = ~N185;
  assign N249 = ~N190;
  assign N250 = ~N195;
  assign N251 = ~N200;
  assign N252 = ~N205;
  assign N253 = ~N210;
  assign N254 = ~N215;
  assign N255 = ~N223;

  always @(posedge clk_i) begin
    if(N224) begin
      data_o_15_sv2v_reg <= r_n_0__15_;
      data_o_14_sv2v_reg <= r_n_0__14_;
      data_o_13_sv2v_reg <= r_n_0__13_;
      data_o_12_sv2v_reg <= r_n_0__12_;
      data_o_11_sv2v_reg <= r_n_0__11_;
      data_o_10_sv2v_reg <= r_n_0__10_;
      data_o_9_sv2v_reg <= r_n_0__9_;
      data_o_8_sv2v_reg <= r_n_0__8_;
      data_o_7_sv2v_reg <= r_n_0__7_;
      data_o_6_sv2v_reg <= r_n_0__6_;
      data_o_5_sv2v_reg <= r_n_0__5_;
      data_o_4_sv2v_reg <= r_n_0__4_;
      data_o_3_sv2v_reg <= r_n_0__3_;
      data_o_2_sv2v_reg <= r_n_0__2_;
      data_o_1_sv2v_reg <= r_n_0__1_;
      data_o_0_sv2v_reg <= r_n_0__0_;
    end 
    if(N225) begin
      r_1__15__sv2v_reg <= r_n_1__15_;
      r_1__14__sv2v_reg <= r_n_1__14_;
      r_1__13__sv2v_reg <= r_n_1__13_;
      r_1__12__sv2v_reg <= r_n_1__12_;
      r_1__11__sv2v_reg <= r_n_1__11_;
      r_1__10__sv2v_reg <= r_n_1__10_;
      r_1__9__sv2v_reg <= r_n_1__9_;
      r_1__8__sv2v_reg <= r_n_1__8_;
      r_1__7__sv2v_reg <= r_n_1__7_;
      r_1__6__sv2v_reg <= r_n_1__6_;
      r_1__5__sv2v_reg <= r_n_1__5_;
      r_1__4__sv2v_reg <= r_n_1__4_;
      r_1__3__sv2v_reg <= r_n_1__3_;
      r_1__2__sv2v_reg <= r_n_1__2_;
      r_1__1__sv2v_reg <= r_n_1__1_;
      r_1__0__sv2v_reg <= r_n_1__0_;
    end 
    if(N226) begin
      r_2__15__sv2v_reg <= r_n_2__15_;
      r_2__14__sv2v_reg <= r_n_2__14_;
      r_2__13__sv2v_reg <= r_n_2__13_;
      r_2__12__sv2v_reg <= r_n_2__12_;
      r_2__11__sv2v_reg <= r_n_2__11_;
      r_2__10__sv2v_reg <= r_n_2__10_;
      r_2__9__sv2v_reg <= r_n_2__9_;
      r_2__8__sv2v_reg <= r_n_2__8_;
      r_2__7__sv2v_reg <= r_n_2__7_;
      r_2__6__sv2v_reg <= r_n_2__6_;
      r_2__5__sv2v_reg <= r_n_2__5_;
      r_2__4__sv2v_reg <= r_n_2__4_;
      r_2__3__sv2v_reg <= r_n_2__3_;
      r_2__2__sv2v_reg <= r_n_2__2_;
      r_2__1__sv2v_reg <= r_n_2__1_;
      r_2__0__sv2v_reg <= r_n_2__0_;
    end 
    if(N227) begin
      r_3__15__sv2v_reg <= r_n_3__15_;
      r_3__14__sv2v_reg <= r_n_3__14_;
      r_3__13__sv2v_reg <= r_n_3__13_;
      r_3__12__sv2v_reg <= r_n_3__12_;
      r_3__11__sv2v_reg <= r_n_3__11_;
      r_3__10__sv2v_reg <= r_n_3__10_;
      r_3__9__sv2v_reg <= r_n_3__9_;
      r_3__8__sv2v_reg <= r_n_3__8_;
      r_3__7__sv2v_reg <= r_n_3__7_;
      r_3__6__sv2v_reg <= r_n_3__6_;
      r_3__5__sv2v_reg <= r_n_3__5_;
      r_3__4__sv2v_reg <= r_n_3__4_;
      r_3__3__sv2v_reg <= r_n_3__3_;
      r_3__2__sv2v_reg <= r_n_3__2_;
      r_3__1__sv2v_reg <= r_n_3__1_;
      r_3__0__sv2v_reg <= r_n_3__0_;
    end 
    if(N228) begin
      r_4__15__sv2v_reg <= r_n_4__15_;
      r_4__14__sv2v_reg <= r_n_4__14_;
      r_4__13__sv2v_reg <= r_n_4__13_;
      r_4__12__sv2v_reg <= r_n_4__12_;
      r_4__11__sv2v_reg <= r_n_4__11_;
      r_4__10__sv2v_reg <= r_n_4__10_;
      r_4__9__sv2v_reg <= r_n_4__9_;
      r_4__8__sv2v_reg <= r_n_4__8_;
      r_4__7__sv2v_reg <= r_n_4__7_;
      r_4__6__sv2v_reg <= r_n_4__6_;
      r_4__5__sv2v_reg <= r_n_4__5_;
      r_4__4__sv2v_reg <= r_n_4__4_;
      r_4__3__sv2v_reg <= r_n_4__3_;
      r_4__2__sv2v_reg <= r_n_4__2_;
      r_4__1__sv2v_reg <= r_n_4__1_;
      r_4__0__sv2v_reg <= r_n_4__0_;
    end 
    if(N229) begin
      r_5__15__sv2v_reg <= r_n_5__15_;
      r_5__14__sv2v_reg <= r_n_5__14_;
      r_5__13__sv2v_reg <= r_n_5__13_;
      r_5__12__sv2v_reg <= r_n_5__12_;
      r_5__11__sv2v_reg <= r_n_5__11_;
      r_5__10__sv2v_reg <= r_n_5__10_;
      r_5__9__sv2v_reg <= r_n_5__9_;
      r_5__8__sv2v_reg <= r_n_5__8_;
      r_5__7__sv2v_reg <= r_n_5__7_;
      r_5__6__sv2v_reg <= r_n_5__6_;
      r_5__5__sv2v_reg <= r_n_5__5_;
      r_5__4__sv2v_reg <= r_n_5__4_;
      r_5__3__sv2v_reg <= r_n_5__3_;
      r_5__2__sv2v_reg <= r_n_5__2_;
      r_5__1__sv2v_reg <= r_n_5__1_;
      r_5__0__sv2v_reg <= r_n_5__0_;
    end 
    if(N230) begin
      r_6__15__sv2v_reg <= r_n_6__15_;
      r_6__14__sv2v_reg <= r_n_6__14_;
      r_6__13__sv2v_reg <= r_n_6__13_;
      r_6__12__sv2v_reg <= r_n_6__12_;
      r_6__11__sv2v_reg <= r_n_6__11_;
      r_6__10__sv2v_reg <= r_n_6__10_;
      r_6__9__sv2v_reg <= r_n_6__9_;
      r_6__8__sv2v_reg <= r_n_6__8_;
      r_6__7__sv2v_reg <= r_n_6__7_;
      r_6__6__sv2v_reg <= r_n_6__6_;
      r_6__5__sv2v_reg <= r_n_6__5_;
      r_6__4__sv2v_reg <= r_n_6__4_;
      r_6__3__sv2v_reg <= r_n_6__3_;
      r_6__2__sv2v_reg <= r_n_6__2_;
      r_6__1__sv2v_reg <= r_n_6__1_;
      r_6__0__sv2v_reg <= r_n_6__0_;
    end 
    if(N231) begin
      r_7__15__sv2v_reg <= r_n_7__15_;
      r_7__14__sv2v_reg <= r_n_7__14_;
      r_7__13__sv2v_reg <= r_n_7__13_;
      r_7__12__sv2v_reg <= r_n_7__12_;
      r_7__11__sv2v_reg <= r_n_7__11_;
      r_7__10__sv2v_reg <= r_n_7__10_;
      r_7__9__sv2v_reg <= r_n_7__9_;
      r_7__8__sv2v_reg <= r_n_7__8_;
      r_7__7__sv2v_reg <= r_n_7__7_;
      r_7__6__sv2v_reg <= r_n_7__6_;
      r_7__5__sv2v_reg <= r_n_7__5_;
      r_7__4__sv2v_reg <= r_n_7__4_;
      r_7__3__sv2v_reg <= r_n_7__3_;
      r_7__2__sv2v_reg <= r_n_7__2_;
      r_7__1__sv2v_reg <= r_n_7__1_;
      r_7__0__sv2v_reg <= r_n_7__0_;
    end 
    if(N232) begin
      r_8__15__sv2v_reg <= r_n_8__15_;
      r_8__14__sv2v_reg <= r_n_8__14_;
      r_8__13__sv2v_reg <= r_n_8__13_;
      r_8__12__sv2v_reg <= r_n_8__12_;
      r_8__11__sv2v_reg <= r_n_8__11_;
      r_8__10__sv2v_reg <= r_n_8__10_;
      r_8__9__sv2v_reg <= r_n_8__9_;
      r_8__8__sv2v_reg <= r_n_8__8_;
      r_8__7__sv2v_reg <= r_n_8__7_;
      r_8__6__sv2v_reg <= r_n_8__6_;
      r_8__5__sv2v_reg <= r_n_8__5_;
      r_8__4__sv2v_reg <= r_n_8__4_;
      r_8__3__sv2v_reg <= r_n_8__3_;
      r_8__2__sv2v_reg <= r_n_8__2_;
      r_8__1__sv2v_reg <= r_n_8__1_;
      r_8__0__sv2v_reg <= r_n_8__0_;
    end 
    if(N233) begin
      r_9__15__sv2v_reg <= r_n_9__15_;
      r_9__14__sv2v_reg <= r_n_9__14_;
      r_9__13__sv2v_reg <= r_n_9__13_;
      r_9__12__sv2v_reg <= r_n_9__12_;
      r_9__11__sv2v_reg <= r_n_9__11_;
      r_9__10__sv2v_reg <= r_n_9__10_;
      r_9__9__sv2v_reg <= r_n_9__9_;
      r_9__8__sv2v_reg <= r_n_9__8_;
      r_9__7__sv2v_reg <= r_n_9__7_;
      r_9__6__sv2v_reg <= r_n_9__6_;
      r_9__5__sv2v_reg <= r_n_9__5_;
      r_9__4__sv2v_reg <= r_n_9__4_;
      r_9__3__sv2v_reg <= r_n_9__3_;
      r_9__2__sv2v_reg <= r_n_9__2_;
      r_9__1__sv2v_reg <= r_n_9__1_;
      r_9__0__sv2v_reg <= r_n_9__0_;
    end 
    if(N234) begin
      r_10__15__sv2v_reg <= r_n_10__15_;
      r_10__14__sv2v_reg <= r_n_10__14_;
      r_10__13__sv2v_reg <= r_n_10__13_;
      r_10__12__sv2v_reg <= r_n_10__12_;
      r_10__11__sv2v_reg <= r_n_10__11_;
      r_10__10__sv2v_reg <= r_n_10__10_;
      r_10__9__sv2v_reg <= r_n_10__9_;
      r_10__8__sv2v_reg <= r_n_10__8_;
      r_10__7__sv2v_reg <= r_n_10__7_;
      r_10__6__sv2v_reg <= r_n_10__6_;
      r_10__5__sv2v_reg <= r_n_10__5_;
      r_10__4__sv2v_reg <= r_n_10__4_;
      r_10__3__sv2v_reg <= r_n_10__3_;
      r_10__2__sv2v_reg <= r_n_10__2_;
      r_10__1__sv2v_reg <= r_n_10__1_;
      r_10__0__sv2v_reg <= r_n_10__0_;
    end 
    if(N235) begin
      r_11__15__sv2v_reg <= r_n_11__15_;
      r_11__14__sv2v_reg <= r_n_11__14_;
      r_11__13__sv2v_reg <= r_n_11__13_;
      r_11__12__sv2v_reg <= r_n_11__12_;
      r_11__11__sv2v_reg <= r_n_11__11_;
      r_11__10__sv2v_reg <= r_n_11__10_;
      r_11__9__sv2v_reg <= r_n_11__9_;
      r_11__8__sv2v_reg <= r_n_11__8_;
      r_11__7__sv2v_reg <= r_n_11__7_;
      r_11__6__sv2v_reg <= r_n_11__6_;
      r_11__5__sv2v_reg <= r_n_11__5_;
      r_11__4__sv2v_reg <= r_n_11__4_;
      r_11__3__sv2v_reg <= r_n_11__3_;
      r_11__2__sv2v_reg <= r_n_11__2_;
      r_11__1__sv2v_reg <= r_n_11__1_;
      r_11__0__sv2v_reg <= r_n_11__0_;
    end 
    if(N236) begin
      r_12__15__sv2v_reg <= r_n_12__15_;
      r_12__14__sv2v_reg <= r_n_12__14_;
      r_12__13__sv2v_reg <= r_n_12__13_;
      r_12__12__sv2v_reg <= r_n_12__12_;
      r_12__11__sv2v_reg <= r_n_12__11_;
      r_12__10__sv2v_reg <= r_n_12__10_;
      r_12__9__sv2v_reg <= r_n_12__9_;
      r_12__8__sv2v_reg <= r_n_12__8_;
      r_12__7__sv2v_reg <= r_n_12__7_;
      r_12__6__sv2v_reg <= r_n_12__6_;
      r_12__5__sv2v_reg <= r_n_12__5_;
      r_12__4__sv2v_reg <= r_n_12__4_;
      r_12__3__sv2v_reg <= r_n_12__3_;
      r_12__2__sv2v_reg <= r_n_12__2_;
      r_12__1__sv2v_reg <= r_n_12__1_;
      r_12__0__sv2v_reg <= r_n_12__0_;
    end 
    if(N237) begin
      r_13__15__sv2v_reg <= r_n_13__15_;
      r_13__14__sv2v_reg <= r_n_13__14_;
      r_13__13__sv2v_reg <= r_n_13__13_;
      r_13__12__sv2v_reg <= r_n_13__12_;
      r_13__11__sv2v_reg <= r_n_13__11_;
      r_13__10__sv2v_reg <= r_n_13__10_;
      r_13__9__sv2v_reg <= r_n_13__9_;
      r_13__8__sv2v_reg <= r_n_13__8_;
      r_13__7__sv2v_reg <= r_n_13__7_;
      r_13__6__sv2v_reg <= r_n_13__6_;
      r_13__5__sv2v_reg <= r_n_13__5_;
      r_13__4__sv2v_reg <= r_n_13__4_;
      r_13__3__sv2v_reg <= r_n_13__3_;
      r_13__2__sv2v_reg <= r_n_13__2_;
      r_13__1__sv2v_reg <= r_n_13__1_;
      r_13__0__sv2v_reg <= r_n_13__0_;
    end 
    if(N238) begin
      r_14__15__sv2v_reg <= r_n_14__15_;
      r_14__14__sv2v_reg <= r_n_14__14_;
      r_14__13__sv2v_reg <= r_n_14__13_;
      r_14__12__sv2v_reg <= r_n_14__12_;
      r_14__11__sv2v_reg <= r_n_14__11_;
      r_14__10__sv2v_reg <= r_n_14__10_;
      r_14__9__sv2v_reg <= r_n_14__9_;
      r_14__8__sv2v_reg <= r_n_14__8_;
      r_14__7__sv2v_reg <= r_n_14__7_;
      r_14__6__sv2v_reg <= r_n_14__6_;
      r_14__5__sv2v_reg <= r_n_14__5_;
      r_14__4__sv2v_reg <= r_n_14__4_;
      r_14__3__sv2v_reg <= r_n_14__3_;
      r_14__2__sv2v_reg <= r_n_14__2_;
      r_14__1__sv2v_reg <= r_n_14__1_;
      r_14__0__sv2v_reg <= r_n_14__0_;
    end 
    if(N239) begin
      r_15__15__sv2v_reg <= r_n_15__15_;
      r_15__14__sv2v_reg <= r_n_15__14_;
      r_15__13__sv2v_reg <= r_n_15__13_;
      r_15__12__sv2v_reg <= r_n_15__12_;
      r_15__11__sv2v_reg <= r_n_15__11_;
      r_15__10__sv2v_reg <= r_n_15__10_;
      r_15__9__sv2v_reg <= r_n_15__9_;
      r_15__8__sv2v_reg <= r_n_15__8_;
      r_15__7__sv2v_reg <= r_n_15__7_;
      r_15__6__sv2v_reg <= r_n_15__6_;
      r_15__5__sv2v_reg <= r_n_15__5_;
      r_15__4__sv2v_reg <= r_n_15__4_;
      r_15__3__sv2v_reg <= r_n_15__3_;
      r_15__2__sv2v_reg <= r_n_15__2_;
      r_15__1__sv2v_reg <= r_n_15__1_;
      r_15__0__sv2v_reg <= r_n_15__0_;
    end 
    if(N240) begin
      r_16__15__sv2v_reg <= r_n_16__15_;
      r_16__14__sv2v_reg <= r_n_16__14_;
      r_16__13__sv2v_reg <= r_n_16__13_;
      r_16__12__sv2v_reg <= r_n_16__12_;
      r_16__11__sv2v_reg <= r_n_16__11_;
      r_16__10__sv2v_reg <= r_n_16__10_;
      r_16__9__sv2v_reg <= r_n_16__9_;
      r_16__8__sv2v_reg <= r_n_16__8_;
      r_16__7__sv2v_reg <= r_n_16__7_;
      r_16__6__sv2v_reg <= r_n_16__6_;
      r_16__5__sv2v_reg <= r_n_16__5_;
      r_16__4__sv2v_reg <= r_n_16__4_;
      r_16__3__sv2v_reg <= r_n_16__3_;
      r_16__2__sv2v_reg <= r_n_16__2_;
      r_16__1__sv2v_reg <= r_n_16__1_;
      r_16__0__sv2v_reg <= r_n_16__0_;
    end 
    if(N241) begin
      r_17__15__sv2v_reg <= r_n_17__15_;
      r_17__14__sv2v_reg <= r_n_17__14_;
      r_17__13__sv2v_reg <= r_n_17__13_;
      r_17__12__sv2v_reg <= r_n_17__12_;
      r_17__11__sv2v_reg <= r_n_17__11_;
      r_17__10__sv2v_reg <= r_n_17__10_;
      r_17__9__sv2v_reg <= r_n_17__9_;
      r_17__8__sv2v_reg <= r_n_17__8_;
      r_17__7__sv2v_reg <= r_n_17__7_;
      r_17__6__sv2v_reg <= r_n_17__6_;
      r_17__5__sv2v_reg <= r_n_17__5_;
      r_17__4__sv2v_reg <= r_n_17__4_;
      r_17__3__sv2v_reg <= r_n_17__3_;
      r_17__2__sv2v_reg <= r_n_17__2_;
      r_17__1__sv2v_reg <= r_n_17__1_;
      r_17__0__sv2v_reg <= r_n_17__0_;
    end 
    if(N242) begin
      r_18__15__sv2v_reg <= r_n_18__15_;
      r_18__14__sv2v_reg <= r_n_18__14_;
      r_18__13__sv2v_reg <= r_n_18__13_;
      r_18__12__sv2v_reg <= r_n_18__12_;
      r_18__11__sv2v_reg <= r_n_18__11_;
      r_18__10__sv2v_reg <= r_n_18__10_;
      r_18__9__sv2v_reg <= r_n_18__9_;
      r_18__8__sv2v_reg <= r_n_18__8_;
      r_18__7__sv2v_reg <= r_n_18__7_;
      r_18__6__sv2v_reg <= r_n_18__6_;
      r_18__5__sv2v_reg <= r_n_18__5_;
      r_18__4__sv2v_reg <= r_n_18__4_;
      r_18__3__sv2v_reg <= r_n_18__3_;
      r_18__2__sv2v_reg <= r_n_18__2_;
      r_18__1__sv2v_reg <= r_n_18__1_;
      r_18__0__sv2v_reg <= r_n_18__0_;
    end 
    if(N243) begin
      r_19__15__sv2v_reg <= r_n_19__15_;
      r_19__14__sv2v_reg <= r_n_19__14_;
      r_19__13__sv2v_reg <= r_n_19__13_;
      r_19__12__sv2v_reg <= r_n_19__12_;
      r_19__11__sv2v_reg <= r_n_19__11_;
      r_19__10__sv2v_reg <= r_n_19__10_;
      r_19__9__sv2v_reg <= r_n_19__9_;
      r_19__8__sv2v_reg <= r_n_19__8_;
      r_19__7__sv2v_reg <= r_n_19__7_;
      r_19__6__sv2v_reg <= r_n_19__6_;
      r_19__5__sv2v_reg <= r_n_19__5_;
      r_19__4__sv2v_reg <= r_n_19__4_;
      r_19__3__sv2v_reg <= r_n_19__3_;
      r_19__2__sv2v_reg <= r_n_19__2_;
      r_19__1__sv2v_reg <= r_n_19__1_;
      r_19__0__sv2v_reg <= r_n_19__0_;
    end 
    if(N244) begin
      r_20__15__sv2v_reg <= r_n_20__15_;
      r_20__14__sv2v_reg <= r_n_20__14_;
      r_20__13__sv2v_reg <= r_n_20__13_;
      r_20__12__sv2v_reg <= r_n_20__12_;
      r_20__11__sv2v_reg <= r_n_20__11_;
      r_20__10__sv2v_reg <= r_n_20__10_;
      r_20__9__sv2v_reg <= r_n_20__9_;
      r_20__8__sv2v_reg <= r_n_20__8_;
      r_20__7__sv2v_reg <= r_n_20__7_;
      r_20__6__sv2v_reg <= r_n_20__6_;
      r_20__5__sv2v_reg <= r_n_20__5_;
      r_20__4__sv2v_reg <= r_n_20__4_;
      r_20__3__sv2v_reg <= r_n_20__3_;
      r_20__2__sv2v_reg <= r_n_20__2_;
      r_20__1__sv2v_reg <= r_n_20__1_;
      r_20__0__sv2v_reg <= r_n_20__0_;
    end 
    if(N245) begin
      r_21__15__sv2v_reg <= r_n_21__15_;
      r_21__14__sv2v_reg <= r_n_21__14_;
      r_21__13__sv2v_reg <= r_n_21__13_;
      r_21__12__sv2v_reg <= r_n_21__12_;
      r_21__11__sv2v_reg <= r_n_21__11_;
      r_21__10__sv2v_reg <= r_n_21__10_;
      r_21__9__sv2v_reg <= r_n_21__9_;
      r_21__8__sv2v_reg <= r_n_21__8_;
      r_21__7__sv2v_reg <= r_n_21__7_;
      r_21__6__sv2v_reg <= r_n_21__6_;
      r_21__5__sv2v_reg <= r_n_21__5_;
      r_21__4__sv2v_reg <= r_n_21__4_;
      r_21__3__sv2v_reg <= r_n_21__3_;
      r_21__2__sv2v_reg <= r_n_21__2_;
      r_21__1__sv2v_reg <= r_n_21__1_;
      r_21__0__sv2v_reg <= r_n_21__0_;
    end 
    if(N246) begin
      r_22__15__sv2v_reg <= r_n_22__15_;
      r_22__14__sv2v_reg <= r_n_22__14_;
      r_22__13__sv2v_reg <= r_n_22__13_;
      r_22__12__sv2v_reg <= r_n_22__12_;
      r_22__11__sv2v_reg <= r_n_22__11_;
      r_22__10__sv2v_reg <= r_n_22__10_;
      r_22__9__sv2v_reg <= r_n_22__9_;
      r_22__8__sv2v_reg <= r_n_22__8_;
      r_22__7__sv2v_reg <= r_n_22__7_;
      r_22__6__sv2v_reg <= r_n_22__6_;
      r_22__5__sv2v_reg <= r_n_22__5_;
      r_22__4__sv2v_reg <= r_n_22__4_;
      r_22__3__sv2v_reg <= r_n_22__3_;
      r_22__2__sv2v_reg <= r_n_22__2_;
      r_22__1__sv2v_reg <= r_n_22__1_;
      r_22__0__sv2v_reg <= r_n_22__0_;
    end 
    if(N247) begin
      r_23__15__sv2v_reg <= r_n_23__15_;
      r_23__14__sv2v_reg <= r_n_23__14_;
      r_23__13__sv2v_reg <= r_n_23__13_;
      r_23__12__sv2v_reg <= r_n_23__12_;
      r_23__11__sv2v_reg <= r_n_23__11_;
      r_23__10__sv2v_reg <= r_n_23__10_;
      r_23__9__sv2v_reg <= r_n_23__9_;
      r_23__8__sv2v_reg <= r_n_23__8_;
      r_23__7__sv2v_reg <= r_n_23__7_;
      r_23__6__sv2v_reg <= r_n_23__6_;
      r_23__5__sv2v_reg <= r_n_23__5_;
      r_23__4__sv2v_reg <= r_n_23__4_;
      r_23__3__sv2v_reg <= r_n_23__3_;
      r_23__2__sv2v_reg <= r_n_23__2_;
      r_23__1__sv2v_reg <= r_n_23__1_;
      r_23__0__sv2v_reg <= r_n_23__0_;
    end 
    if(N248) begin
      r_24__15__sv2v_reg <= r_n_24__15_;
      r_24__14__sv2v_reg <= r_n_24__14_;
      r_24__13__sv2v_reg <= r_n_24__13_;
      r_24__12__sv2v_reg <= r_n_24__12_;
      r_24__11__sv2v_reg <= r_n_24__11_;
      r_24__10__sv2v_reg <= r_n_24__10_;
      r_24__9__sv2v_reg <= r_n_24__9_;
      r_24__8__sv2v_reg <= r_n_24__8_;
      r_24__7__sv2v_reg <= r_n_24__7_;
      r_24__6__sv2v_reg <= r_n_24__6_;
      r_24__5__sv2v_reg <= r_n_24__5_;
      r_24__4__sv2v_reg <= r_n_24__4_;
      r_24__3__sv2v_reg <= r_n_24__3_;
      r_24__2__sv2v_reg <= r_n_24__2_;
      r_24__1__sv2v_reg <= r_n_24__1_;
      r_24__0__sv2v_reg <= r_n_24__0_;
    end 
    if(N249) begin
      r_25__15__sv2v_reg <= r_n_25__15_;
      r_25__14__sv2v_reg <= r_n_25__14_;
      r_25__13__sv2v_reg <= r_n_25__13_;
      r_25__12__sv2v_reg <= r_n_25__12_;
      r_25__11__sv2v_reg <= r_n_25__11_;
      r_25__10__sv2v_reg <= r_n_25__10_;
      r_25__9__sv2v_reg <= r_n_25__9_;
      r_25__8__sv2v_reg <= r_n_25__8_;
      r_25__7__sv2v_reg <= r_n_25__7_;
      r_25__6__sv2v_reg <= r_n_25__6_;
      r_25__5__sv2v_reg <= r_n_25__5_;
      r_25__4__sv2v_reg <= r_n_25__4_;
      r_25__3__sv2v_reg <= r_n_25__3_;
      r_25__2__sv2v_reg <= r_n_25__2_;
      r_25__1__sv2v_reg <= r_n_25__1_;
      r_25__0__sv2v_reg <= r_n_25__0_;
    end 
    if(N250) begin
      r_26__15__sv2v_reg <= r_n_26__15_;
      r_26__14__sv2v_reg <= r_n_26__14_;
      r_26__13__sv2v_reg <= r_n_26__13_;
      r_26__12__sv2v_reg <= r_n_26__12_;
      r_26__11__sv2v_reg <= r_n_26__11_;
      r_26__10__sv2v_reg <= r_n_26__10_;
      r_26__9__sv2v_reg <= r_n_26__9_;
      r_26__8__sv2v_reg <= r_n_26__8_;
      r_26__7__sv2v_reg <= r_n_26__7_;
      r_26__6__sv2v_reg <= r_n_26__6_;
      r_26__5__sv2v_reg <= r_n_26__5_;
      r_26__4__sv2v_reg <= r_n_26__4_;
      r_26__3__sv2v_reg <= r_n_26__3_;
      r_26__2__sv2v_reg <= r_n_26__2_;
      r_26__1__sv2v_reg <= r_n_26__1_;
      r_26__0__sv2v_reg <= r_n_26__0_;
    end 
    if(N251) begin
      r_27__15__sv2v_reg <= r_n_27__15_;
      r_27__14__sv2v_reg <= r_n_27__14_;
      r_27__13__sv2v_reg <= r_n_27__13_;
      r_27__12__sv2v_reg <= r_n_27__12_;
      r_27__11__sv2v_reg <= r_n_27__11_;
      r_27__10__sv2v_reg <= r_n_27__10_;
      r_27__9__sv2v_reg <= r_n_27__9_;
      r_27__8__sv2v_reg <= r_n_27__8_;
      r_27__7__sv2v_reg <= r_n_27__7_;
      r_27__6__sv2v_reg <= r_n_27__6_;
      r_27__5__sv2v_reg <= r_n_27__5_;
      r_27__4__sv2v_reg <= r_n_27__4_;
      r_27__3__sv2v_reg <= r_n_27__3_;
      r_27__2__sv2v_reg <= r_n_27__2_;
      r_27__1__sv2v_reg <= r_n_27__1_;
      r_27__0__sv2v_reg <= r_n_27__0_;
    end 
    if(N252) begin
      r_28__15__sv2v_reg <= r_n_28__15_;
      r_28__14__sv2v_reg <= r_n_28__14_;
      r_28__13__sv2v_reg <= r_n_28__13_;
      r_28__12__sv2v_reg <= r_n_28__12_;
      r_28__11__sv2v_reg <= r_n_28__11_;
      r_28__10__sv2v_reg <= r_n_28__10_;
      r_28__9__sv2v_reg <= r_n_28__9_;
      r_28__8__sv2v_reg <= r_n_28__8_;
      r_28__7__sv2v_reg <= r_n_28__7_;
      r_28__6__sv2v_reg <= r_n_28__6_;
      r_28__5__sv2v_reg <= r_n_28__5_;
      r_28__4__sv2v_reg <= r_n_28__4_;
      r_28__3__sv2v_reg <= r_n_28__3_;
      r_28__2__sv2v_reg <= r_n_28__2_;
      r_28__1__sv2v_reg <= r_n_28__1_;
      r_28__0__sv2v_reg <= r_n_28__0_;
    end 
    if(N253) begin
      r_29__15__sv2v_reg <= r_n_29__15_;
      r_29__14__sv2v_reg <= r_n_29__14_;
      r_29__13__sv2v_reg <= r_n_29__13_;
      r_29__12__sv2v_reg <= r_n_29__12_;
      r_29__11__sv2v_reg <= r_n_29__11_;
      r_29__10__sv2v_reg <= r_n_29__10_;
      r_29__9__sv2v_reg <= r_n_29__9_;
      r_29__8__sv2v_reg <= r_n_29__8_;
      r_29__7__sv2v_reg <= r_n_29__7_;
      r_29__6__sv2v_reg <= r_n_29__6_;
      r_29__5__sv2v_reg <= r_n_29__5_;
      r_29__4__sv2v_reg <= r_n_29__4_;
      r_29__3__sv2v_reg <= r_n_29__3_;
      r_29__2__sv2v_reg <= r_n_29__2_;
      r_29__1__sv2v_reg <= r_n_29__1_;
      r_29__0__sv2v_reg <= r_n_29__0_;
    end 
    if(N254) begin
      r_30__15__sv2v_reg <= r_n_30__15_;
      r_30__14__sv2v_reg <= r_n_30__14_;
      r_30__13__sv2v_reg <= r_n_30__13_;
      r_30__12__sv2v_reg <= r_n_30__12_;
      r_30__11__sv2v_reg <= r_n_30__11_;
      r_30__10__sv2v_reg <= r_n_30__10_;
      r_30__9__sv2v_reg <= r_n_30__9_;
      r_30__8__sv2v_reg <= r_n_30__8_;
      r_30__7__sv2v_reg <= r_n_30__7_;
      r_30__6__sv2v_reg <= r_n_30__6_;
      r_30__5__sv2v_reg <= r_n_30__5_;
      r_30__4__sv2v_reg <= r_n_30__4_;
      r_30__3__sv2v_reg <= r_n_30__3_;
      r_30__2__sv2v_reg <= r_n_30__2_;
      r_30__1__sv2v_reg <= r_n_30__1_;
      r_30__0__sv2v_reg <= r_n_30__0_;
    end 
    if(N219) begin
      r_31__15__sv2v_reg <= 1'b0;
      r_31__14__sv2v_reg <= 1'b0;
      r_31__13__sv2v_reg <= 1'b0;
      r_31__12__sv2v_reg <= 1'b0;
      r_31__11__sv2v_reg <= 1'b0;
      r_31__10__sv2v_reg <= 1'b0;
      r_31__9__sv2v_reg <= 1'b0;
      r_31__8__sv2v_reg <= 1'b0;
      r_31__7__sv2v_reg <= 1'b0;
      r_31__6__sv2v_reg <= 1'b0;
      r_31__5__sv2v_reg <= 1'b0;
      r_31__4__sv2v_reg <= 1'b0;
      r_31__3__sv2v_reg <= 1'b0;
      r_31__2__sv2v_reg <= 1'b0;
      r_31__1__sv2v_reg <= 1'b0;
      r_31__0__sv2v_reg <= 1'b0;
    end else if(N255) begin
      r_31__15__sv2v_reg <= data_i[15];
      r_31__14__sv2v_reg <= data_i[14];
      r_31__13__sv2v_reg <= data_i[13];
      r_31__12__sv2v_reg <= data_i[12];
      r_31__11__sv2v_reg <= data_i[11];
      r_31__10__sv2v_reg <= data_i[10];
      r_31__9__sv2v_reg <= data_i[9];
      r_31__8__sv2v_reg <= data_i[8];
      r_31__7__sv2v_reg <= data_i[7];
      r_31__6__sv2v_reg <= data_i[6];
      r_31__5__sv2v_reg <= data_i[5];
      r_31__4__sv2v_reg <= data_i[4];
      r_31__3__sv2v_reg <= data_i[3];
      r_31__2__sv2v_reg <= data_i[2];
      r_31__1__sv2v_reg <= data_i[1];
      r_31__0__sv2v_reg <= data_i[0];
    end 
  end


endmodule

