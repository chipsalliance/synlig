module dut (input a, output b);
	assign b = $unsigned(a);
endmodule
